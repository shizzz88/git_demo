��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"If�Q�L��A��l�rX��1�򕑘�����G󍹭�!�V1���B��?ھ����)DG��󀼶��D-�Ɠx��;�y���z~�F����0S��>v��᷼-�xiq���I�Q͊DK^�'���xW�(�h�����E�<�6z+w}�`uz�ީ���tP��vO�(��C�!�������v���w��{��[�]���,}�(Fr��;z�ȐT+
)M9�'���@���|���-A�â%�`����<� -�.�b������N��|�8t=/1������m4(jP�`�{��L�Z[�Q��D�9���!�сJ��h��6������In���t��F��D襴X�,q2Y6x�T��T9���|b���K�k�j�P��A��2�%I�������<f�d�N3l�V���QѠ�a�V�����m]����T�S0���Cү0^�J!V|!M�T����f�L��p��g͟�TA�Hx�l�B�k�ԋrf �;�#6� �6��f3-3� }ҚZ��E����Y�U3`@0� ���7e�7�d�G꛷�v�ل�6�a�����{
��!-g�l�@WG�-Љ �ؾa�{��LU �����(��K�`�S�ݵ���O�O^��tDF�:@�	�����،N�38.b8ے[��P)�Ͳ��3����ЕRe��ԍ[ϱiP%��:*�=$Q����B4�k�PI�.ŵ�O*[��j���)��!x��m>94�a��� �UE-�������A�'�~Py�ྵ��Pj�ߟ��]'���5�������r�m,t;�����^�3d_��n�b���G�ZDa�<4�
�Ee:��b�奜�7�=��1�l��+��`�+\�Ê=�<ǐ�F�9I7a����	�k0П���Z8��AmY�.+��%$g�P�?�������H��a��M�� ����c-����9�$	��u2 0�n��7EXsk�h?��eْ<|�Ѹw���#�+p����C9�5�á�{��q}�}��st����݂6R��¨Gd#�ѷ$Ws���Zѫ�bب�Ч�N�YԞ�mw��E!7���.��3�b���*��~@�6JN8�>K� \&�o��Y<"Є1!�-V�cae�����w��UR{�'���#�c�:?+U����������3@��o[���q���D�Y�#�ZBPJ�^������__g�f	���}�>�I�Q��Y:�?V����2��s{����*�s�i"��Fnp�3��_��gi���6K���)� �zN\����-���Yo�x�����.���4��dE`��L���lH�"n�E��Kxm�K׶C{� (��Zw�Yg=|LIU[sc>�X)�,q�P��#�A�$�!�~T4<Z�,iS*����M���q"���4@w#�!|�f�����af]���f�%Ϋt\��A�|���̄��R����į���%7��&�����M��L!�x�K
���x+�-�𑫻�&����(���� ��5������I��(\1���25���H��`Anw��e����Yig��ky.i�
��7&��'x���n�]G�c��E��A5k0��P�'���l�m)V3�Sz3hlV�g�����ұ#��O �v����N���-##�V3D/;�8�H�չ�e�}��a�I*��Ƶ6`��EȋZzE�D+;|E�p1�jX���ɗ��t�$��u��Ω��x�<�k���	�����X�b��&��tI�Oވ���\�Z����� ױ��Q?�Jp$���xp�E ���}3��e�۠�}}���(�Q�O�	Y�������?�+ln���Py���_��O.�%�n��uBE+(�x����Oa��݇�.7q�J��Ȍ�k���20�r����/�A���q	��v�ŏ����rE�l�*ߑ�!��C����aJ�b.�܀y#M�*���}Q�nނwy����=��R�wp� I�`�řz�fz&Cل��A^3q���#���c�`��|�7�;**�|�&=e�/<�D��l)�.>�kJ���B8R*�!
�j�g��$�yTD��r�ҩ��)��m���B��X�򦕱'�9~�5��_7��B%�G�م��d��j;5���73�^�����7�g��!�:��hP�4��߉��#Os�Z�lC�m��Z H4���DS�Ă���Ƥ5�G�����&̶O'S�׉f�L]B�{������#�wg0g���e�"  �my���Du� ;�҈�xI�o�%�A�\A!ڣ����).��v����ۘ�R�TBV>��Ws?���|�5Ӽ9k4�]�0�F,H'S!�fem=^J��0W��C�i����zl+�D;�p�q����m�E����X���A�b�	Lq�݄ġ���Z9,ȋ��%>���a�
-��x�ۉ�-��a P�X�w�l$2��ӫ�Qo{j>�x�-�s%boe%�Y���E�آgG�ƨ�����=�ݰ 5����ԅ����d�p9;֩)6���H���=���X�/pA���0�,��"u?Y�z�6�d�}Bfe��'X�l5�F5�k����f�z�k@��F拴��A2���L�B������u� �sT���L��v?Y� ܜPA���pN��g8j����=`��{9G�������,�1�@()ѡv�"�rG��'|���J�aQs I[���843�8FCU�nD3���� ,R�&7�k�븬��/�v�#�~uXd���%��-8I9D��7B�SF��`�_�ϋ�;Vq�CIg��;�0˲7:C�r`�7=U�#;�JI@�wq���kL��S�կ��ZK��&�#�����Ek[F���u�% �}��t�w#U���<�~�ՈN�N;���������o���gva2��8�(�ؾ�]�E,����lҼ�>�_q��_"���oߘ �о�r��@2Ī��6e�H��j*�������obl��hJK��v2���`�c�΢|R'fZ"�P�2ک@��.�;./�Qy7�|	1C�8���$��r���^�r�)~8��>h���y�Y���ΐq��?7c������@'��쵺�?k���eC�2%�5P��13��)�����,߆�WhBE8��v ��>%����Z�P�����!� ��Uq��L��$V�}8���3�e�l�u=�\�t�ڑ]%Y��(�V���Kw]HB@����=R�J�����2�֌�w���ւ��a{+�:JW)��,�qbΎ��"��A�Aы֘u��[���
��>E!jY0�]�dw�;�
�A������N}�M_�1K�%�d�Z��93�
6/�Ɖi�O�v��%��x�{H�\±�L�������(��y�Pr����~�|d��Q�<hl��d�b]���sl�:��J����*}��ĩ��Z|�N��7��(��+�|�æ�݉/�I�X�w8����>1����B�^ef
�F�)�kYa��Xa�&c��Nx#1տҷ�����5�;Zr��U��� �U��e�Wɏ����m��6�PУ'�_'�ũ��2�^�0w�����s=��wM����ϖK�W�s�]o�I�6f�7*��.�*8!�	��q��/.��� � i5��,��K��Ǥ͐��>4��@��"�zkx��k���2�����TS_�EFpY�G��jml�8ᐉ��lr{"_N6dy��RG�Q�z�:cn'E�5���?�\�KiE�����v���4ĩ�I-����9�w�$���E��_=����Bn�ꮎ�^㘿���y}+'����ͣ��~��B+c���H2����kʯ���_J��ʎ�$}&`|���Q���Uj���ݯ�e�i6�YJ�+��ϥ� O��W�8�ֶ�(��A���Ʈ�0���`^���k��uZ�q\��/�a )��
#�G��EQ/L�O����+Ec�b�
H	�T����Jw3M"��]�%��ܓt���qxmNNL�H����=����|�s���y��j�;0;1r"UvB��� �m>6_�VkfFD�]�텾�z9� ��(qG1���|������I��"�~:t��2�vuc�{m�z��4�᠀KKT- ���HdU�#Fr+�IM��C�&f��:�~�'R�ߥE�]xgiƽ���#m���.dvYT���ޣ	3	vכp�/��\��1��g��c 81
�h\�*pf[| �,J�Ir������ �'���+�)�	��|k���\p
d:}�aC���Y5H���� �S� ��6�K���`K*��*�����Ļ�U�2���Ay�M:��L�zS��ܹ�okD�K�Q"ʹΜ`U�6�[�����6շ���W��2�Od�Υ���Kbp�kx��!�t	�.��+A��#�X��xoѭ ��w��I�Ľ�rV.C��	V�	�^�㳄a����.e�$��>�3�v���3,'��I���׮�����a����o�i�l^��@���E�>��¥H�C���R��n#Gn������P�d��7��d�f'��l-xg�S���B=����9g�h��m6e�E�:HELE�1���{��U�>8w��C��zL��l>@�Șt��r~���� \�MT��0G�ܶ��rG���sl�}j���������ͪ�XN$R1��R��<Wfj�	�N<�ī���ৌ�>&Y5g�4}}��G�b%�*!�,}���P�Y�%����[�+� �F )W[�K,��4��eb�˔�)�Tb��V�Ȁ��m�h�1�<p���)�H_�L�K�̗�^p�Yn���� ����AYD�7��N�|}�������SB�Al2�n�Me�E�-��y����E>��M���(ˌqUQ�^i}��)�Bʻ 1|N�Qī�;��Q~����;�e�������z���+�V��tt��v4�),�}�ԱM4���K�Qt��r? ,��8��n�n����BrE��Z��oO9~ '�������	��;���Ay�cxQ��B�5��x���HQ��\���R�xj(\i�Ngv��C���9�.$0f~+,��{����1�yt�@�b�t�O���>UV`�����D�<$Vq�j'�5��/l�����+;<��TD?PJ<%�[WCh.��Y$ntʮBY!| q�$H��Ϋ���y����e��f�?�<*L�J���C��b��}yY��G�NSQj�o�^D��|i}���q%A��g ��цׂ�I=��ߞ�Uu��LE��v)�|z��DU�R��U�����^H�CzmS:���|^�g�Fb�����V��-��Ubaݢ��(y�)�SD&b�HǦVRz`���Feפ�ǣ��<:��n貸�V�5���T�R0 �7�����Lm��������Q���\��LGȦ!$�3-�1অLo��/��U�`t V��MB'xg�F�:�f���p��wZ
gmż"�!A�EB�p�y����G�ǿ�A)(�1�k�p9m�bQ�i���Y�c
$AK��C��D�Ac�֥u1��X�n_��|��!����\��#MY`=�;�k�<�{{���
�ro_��^NB:,�T���%�#8K�uk��I\>@<"�q��1���lh����Ō��m���'�WR>w@�����k����V� w|!���m�4:���խd�b����.��/�
��>������Qxa?���&�{Agˉa%[ʓJW}���
Z\`~&ҿ}��r �.�$�r�g>w��=wq�g��A=V3�����4�#�;��kҝ��^��Z� �yg��>92�C����-�;�_��+��ց��KN�l�?��m/�m4�?�F�>���16:r��FF�G̵6�l��U�i�,L�jV.v��C�A d�~��R~��܇���^@cb�!�F����/���\ד�Q+����=1ZT���f�}K�~�Uf3+�C�)'��"�Q�a���9q�9,���Qȱ���թN��7��xD��"����&���LvP'Y+r�y]��։;��jū�8�H���F%B�Ҽ#3/C��-0�!_���Ҍ��@ol����ƘW�QN8���}�+%���cj�|QPF�M�-h���0�Ҟ؃�[� Z��嫑}�:�1�4�
�]�,�m�����=��ʿ�ޏ����')�tR�+�H.�f��x+�e�_����_�^�+�K�wb!��S����-~-�7J�.U�h��WV�h�i��q���`<誔-"|�v��
3L�	�(i���_@�\�(��d[-M�C�MK�FX���pV��Wۚ���m;<�I�pb�GG��&�Fh���X��>�W�a�(��/���Z%�P��T�>��:���N�,t�CMin��'߹��"��nJ�ȱ�"�]@r�+F����N�,�{m=�j�	�}3�Q;7 �8vr����~�d�ԧ�+��1��.�NQ��F/<u�%ܥ,Z\X�� �6uD�ۛ��̂�m���� A�{7��(�s ����W�J|�A�'r؜�Ϋ�Q��bm*��jh�����`�"��i�0'�a�GY��ok�OnA�O�>?�K']��{:�͔݋�mx�]��4N�>����Gd��%N��"ΔY�(_&���F�>jYA���]��V��C>��X�]ږ�0�P�Y7�O/3,c���\��N�#W;�����/�C*��p^T�Bp��M�X9m�)h����W�i�
E1;P�-PpP��<e����2�m��1�\�� ��U�U��+�8���M���D���]&����F�4v<mݦ�T�<!CT�Ұ��a�x\Lkߧ���lU���8Z�TR�p��Z0`eRY�����)�����db-��Va��ˮ�?�7�'�.{Ӹ���,bNK>-V	�|��ǡ�$����잀v)H�NU�����+��+�cx��n/[��B�E"W������N�I�-P3~Ochu@�����c���l>�P��&'!x�[��@�2�$�ң���R�h��<3^�؃"��͒ �f�F�z����"ϊ���pUk_�I������'<p3V����%{��VM�Us}����N���,��!j pr�[��]���%ͺ����b `��Pb�Q	s���<|ZNE`_�v�ڍX��&2R7��ä)F��D�s��(�����.f��s�1<V�[�P�	��:�1�y��V�PF�y�f����&�� ��2��h@���]X�0'u���|bt֊-�{b�sk��u��/�G�	g3p58�-������)6s�,)g�Ø���w���8���Z7ɜ��/dn?���:���5nƵ��L��"�O�Z�I��r=�*g�M�	��v�K,jW��@v��"r��9��Y;���͑���=F�_$TdVyC���<�d��'Q WS��U���6�DRz�U���+Ж��X�n�o�:��aw��ԐN�>�5�~�6��VNN��Lbt?^C���;�D��_�R��+�,$q�"��G�ۅD�Ŵ�T,O�^�{l�?�b��$T���k�}1?R��f&�M��bn2��t��ʸz���UY>�val[8]Jq�O�B �1�+^����ޱ�?��z������E�DsCMy���F���2 P�2��+����:Y�}*�X@w���ь��x�Ɂ\K~�T��8$L߀�������項�49M>Moe:��g�=���6�{�o�����?T_�6�����(�¹,G;z�5/�3��?����p�eU�����8��i��Ԡ�:g�X�h�tX4��b�%�'�p@��NF���L���[�9���)�O����[Y�Ղ�)�}Z<U'��63�S�n�%֚Q�ZV�J��b����Z�|`�+F!p���������ky��Z�m�Ė=�.�'���n�tO%�'�s��ld�ND1�����Bԟ�����2�M�Y�o��!2�S�¾+�%*G�ʙ<�Iu��+�/%�JFsv�~yC+p���Ŗ�+vk�a�)_Y� �,N�3H��P�{�V�`t�2� S?������!6���oږ2D1�����ʂ
o�E'N��;���l���Gb�Tx�5x3�G�M�=����u�0K4X���I�h�v�ԁ���QVܔ=�h��.�f�RX��=^#���{	�{[2�T�;��u�OVq�Kb-2Ta'dE��LN�K'oh7\��޷�0�S Ϝ�qi��݂�N�zKȎj+��BH�Q�CFu��h�|��{����*�n?a�7�6�h���	0LƂ#?n�6k%KCWP,@Կ�I>B'mk��>��n�<�,A� �� �{���.D��f��n�i 婙��R�`��:�X��&���c��鴳8Q��WM|'��]���H�8AM�r���g��a:I��\�JlKH&��sN���]�g��
WG� ʞN*�����dX�R|�M�tR(�4�b]3t�T ��m���\<���FGrh�S���9�NpC�����Wǣ��QjO�Y*��g��Na�[�pO�uCiZ<�^b�DQ���|��Un2��u��+�x)e��dO�[|
���&��o����:�Me�KZ��Xډ����}ٛlf΢e(�|Ї�<��=�Y$�Gp�d�Aąt6��e�0�r�e�
�x�̠Y8��W��+S�jݘ+��8�h�I����x���O�RJ�⁗��ӛ��H|��>���h^���Xs��C\��P�� � ݰ�B	l z�x?ư��v8��t��
��L#��R"[6�P;5�(��>`1d=̍S�G�O����D�J����� ܜ>-���Q哨��4�u�ݥ�ˎnM���$�i�P�)���wh?X����|�8��B�w!<��.�7��*Eߋ����j���.���=㽾�ݡ]��͠!�	,#~��5eG,A>���'�V��8h������~'dD6.6��H��F�La���UP����K�T|�f�H������	m>���.'�o��Z���za��H��,�b��]���.s��@��@�����
9��;��.����QH���q�����t���Qbn��,I���E�`��5�T䑘����q`G4D����0��l�}�d�K �|ٙA��Y��|�˘��"�6�Z����&�����	����i;T]"�]moOa�`V��L�¡]������;y�Y �`H�2���O�9T�"���p���M�)��»z�A\g������I'=�rƓ�u�§��E��Q�O������	<{SQS�w��t�/��R)q+c�"������QjUͷĻ�*��VzF�w�B��A�����_S�Qų��5P��%����ES������e/T(z_Bt'Bp���.����mq^��C+��%�W��J3�^�p��]����)}�L�~�2_������_h��P�1$���u7U�$�-,q~���X[d�<��b�Dӏ)����N�Ή$]�I(�m8��F��T�Ɲ	ȋ��~ذ@:y�vA)o?8�����I�������י]�T�R��d��)VV��y��g㥔3���>�ĮF�eF �s )�[}$8����5Só�<I]뽫���B����#��.��I�ĬC�[���y���=���|v5}�JD�"��v��� �>4�~;n�.��dڑ���� ҉H���h�G?u�עG�tP�\Ǜ�uPQ�I�x��8
��9P�{�&�E$��h�1^J���)9��ɓ�Pn�"ȱ=���M����.�
h�_Ga���2\�@PI��.�����'j���K��j#�ח:���^-��K�Y��'k�
ʚm%'C���������#�L6Af呏�erA�'�n&囉��U���`^8��ը\�M�%WE�28��*кs<;<����I��+]�;�#E��^>ԁ �"�ͭl֪�*�bǓNm�??�C�]-��"C^X��nXݯ��=�N�qt�+zj��;�ֻ۔���hs3d��KJڦ�E �]j�վMpZqu�:�;�5���d�G�������)`�w�;���cs���&!.�z"� �<����;�M�>�f���gZ�EgPd' �,�/�|_��g��#U����>�1!9̄�A���䍣�+��nZ9})�[���H ��-�8G�Cu3O=������I�ō�î��5��k�q&��v]�L��Zۛ4��6l^i5���F������&BY�������v�.�cB�4�g{z�
�jۨsZ՛��I:�-����X�B���@�9���Ѓ��	��4��e���B�0�k������{\؅��8���`���YO�l���=ܠK������:�n��6�%�㯂>�;LO��3��f�-+�N�BP�,[8�lI��lR�)p�xx�ti���7��*�8�Ws^��~��/3aJh2��<Y�v{@���+�Os@�	4��F#c]�����l�s��AG�F>�ȑ������[�aL��X���=����a04���9")�;���5��3t�UC����Z8���_�|����`KҘ&ՕD�h�U�x���y5��-�Ԗ�Y� ��Ny��8���$��|�Nr?�x�R�~V�ix&��_����-e��=���n�뙜�0�7�>�a�X,pVI�lD���|�7`�(1q3�)0��İi(�~#p�Zn����r5*9_C�������@l1�L���C�����W���v�&`�<�Xi�S�Mf���>�KA�0���M��r�n&�j�d�a�p����|���k��{�[l[/��H�-@���"��зoH�jr%����}�Ļ#� Hg�cL�@'�&�{��@�(g�`��jt���ePq��L`C&A�N��Y�Ws$¹̬�c?�]�7�9�;�{<7�t�¤�%-3�؇�6��1�7��M\F}v�ګ�N/-��e�1������eOω�h�b����w�5>���^yd�h�"��s���x	N=.1�Co�Z��7b����Եi#�K��rU&8�b�����A�^E��:�g�>O�}<#F��P2�]��}R�>���ٱv�l��&̯�s��F�ܳ�� ��GF5�߳\���y��z�0(�����N*���e�0�ߚ���4�et������h�Ι�:��Z�^䩒�s�����w���ɚ8�zK d���_�����Ъ�Љ���/�=�8���⊄@�{����/�NR�{����g>=�6���9�5Fn��C�����qo���&�ﱻ��
"r5�Bmuý!�6#ĝzr����>+t���<�[��e|��w� ���Bi�zKK�l�$JÞ"k{��1Q������xzU@��8�����1�
��oY���v< �&� �=���2M$�YO*���!G
���Y�L��=�
ȸ��P�~I����@��#��>��i��1����#�v���}ň��CqRldޫX D�zK���@#��I�F��Z#�~7H���8�p`�@O�(�� �+P� �[�jW�D�7�8�Gq}~�c�^"�vrο���-Vԅ��60���IY����҅��Iy>[Ax�@����b�"�{�㈔�~��O�����oH冽	d<o1������'�~�����,޻�?���X(���p�n"�`�b}H��l�\@]�<���P�/�x�!��M��3�v{2�ט�֒���0#�k�v�P�Ж̢���L�K�;��%��Fk�d�<���1��\N�����y�\;��E:xե����薨�	��l�&�F�ɠ�e:�h""�w�[�@a�~�){�aK5�R#�I+��t՘�؁C���TF� ��C�T��\�%Jl ތ�9����m�[������]�G?BY�t��B���@�궥u�Hi1q�;:ٿr�����.�x%U%�ٲ���o��=���]v��p>ѷ;����rC��s�����\̩;�����)��k0M2�P+�c���R��ɠa�l����K|b�C�df�A��=
1�U8Elr!p���˺e�_�	Ut��\��IAu~!���"p�a�o�t�Mm:vVi� yE�'�;t\9�����T�Em��}�����]��/c��㫘f�������K��qsb����>�ٹ��`�Y�A"!~@�L�%����.u|�J)c+�v��d7t��.e����>�-]���j��܆���*AGMdEº �K���h�#r���*#��A�L@��s~�׍�`���O/K4m)�bX�+XJ��hٌ��ë�⁶�Rh�U�\,'�܊�R|����=��l��*�2�H��'d�|��۲L��ơ(�~H��d�9��W#��Zf�T>�u�ҟA8���w�'�q�5h��t��Q��N�0�]��S`П�_� <��xj��-ǚ����͔���JP��+��S0R.�CԶ��pMc��5����B��t4B��t�=�]i����>E��P�u�ߠ��2Q�&����A�� ^S�(�����R4��8��h_�D6Y^X/c73��P}.t�/S�:cP`�\pەo�)�����E~Y�pV4�;C����$����5[ ֝��6I�����7�&�b�Jk���X��7�!����U&O�W�P�`�Ck��*�D��͝@#@ZXUF+Z��0�O��)pj-��4
e���0<"2��kϞ���c1�زf��u��ɠ�w4�ǃoX�����⛾������G0N|�[1�ԉWA�W���w�f�V��Ǎ�P̖V�+�R��E�J0�T���_2��I}��y��C�ȁ��h�5v_/.gZq����p۔��<-���h�����Sd��ƥ_��{kbD5����:�]�Q���V���%Z��\�Fu��P��6����AX)�.p�Z�be;J�AQ���"i�ӟ>���4+-�_ �S�go� ��k���|�*��kau�c�PBK~sP%����-X�D!���J$/'p�T�0����Ol���)t��|�*��e�n������ǲ�T�ew+�0�������&��Z�h�u_�'�Td�¡��!��W�C��irM�!ռ
�k	��Ҧ���?K���
=rq�r�X~��`|�����f ��tP�$PB���[�����>H�'��g��۴�ωr�H?V�L#�*�����>�\�}.#~s�碰����3b�6a�٨?��$-�y���
廌�����3X�/S��"Ʋ O���N�U�ȉc ɳ|�^m���)�Z���	������-���֕�s���ia�D�L��G	܍5�XZ��P�`��oM�3�lT�������ٗz�и�_�.���앇�E��?@�����[���b�C���� }A.�š�F�.x�u�i��1h���\qNW�h��(YB�k�R��!$x����!:[2����b#�y�Z���F*{�6�69�����p���G�rX%���d\lc^�u��h���ȴ� �����5�_�}�G��i�3�5�f�@&L��m���m��WB,7b,mtx?���x���5�+m/�^��Ա�*܎B�)R*�e2��KlGiF�.1��`��U*b%�Cb�c��r�L�4mL��A�^k��0��)��(jfN.��i�7m>���M���w�X�1J�[�Y�!RG�m4?t��np+�gr�^��2��D�S�^�K6��P�R+�\b��G��6�5�T��D=(�wLQHpF@�'�|�x��G������n�	��~�4A��y�[W���(��j#=6~ŦO�1�J�f�L��S
z����e���*�^mUf�|�'�%(HG�Z���>fƒ�:\��Y]��*o���o���5@|��n���/�� =s�<z(���n	����W�VĲ��N�U��7?2�7��D��40�˻�0�B%{��׌e����*�]�J6��J6jF:b���Ѩ�0VL�Qk/���lrA�j]�Xb���JJ�hg}�Է��~1��;���_�ٜ5*�	@��t�`����X5'#|�Y�қ�Ĉ�B2�$��OZ�
��|j���O�K�X���cL�-�mO��P7uG<�P�$b%��
18Ң��rz�[��;'d e'̐�n3Sڤ��\�m�Yq$Ԋ,�FG��k��f��&�=e�z6�b��*��n�����H�����{m4\���=1#7f:��Ѹ� �.�m��(DO���>h_w3~^�B<�\�P_��%h�����?n	~�D�q+��©�b1/�F��ܽ�P"��:����ذ��?�'[�#�=�'�����V��=Z�v���vq�TT���.d���Ө�����٭�������:Zϣ��X!5}�-\aV���x��������
�He��%nc�.٘��ܨ����j�36h����L����#{�=*˨���BM,��5�G�JmlA�' ��9g���������ǡnyl��:�;�,�=5dU�@�x���w�b��Ch�.z�ʋ����R�R�Wnn��rI�+�ѓ&�i����,����AO;�&�M˭�ĺ9�^��!R��A&?�M?�%�2�a����/9'@Y�Ni�ؔ�~C�/��Z��٪T����.tIY�u�D�5F��Mo��*�{Q�dKlQ�u�P.6��\�I��v��[�_3r>�QRCY��&u���84޸}]�eܽ��Z�[ ��g��\��{2)K�:��;&�F�hL�$U��)��#&�i�A��O.�݁�	����*;69�5�|A��h�����6�s
`��f�p���'u��}�ì�E�X���Or��/�x�K�2�+����g�A�@�ٗh�����x��n<��jAc�p	a���P��+Ճiw_cL@�"������0E@�u���Gi_+�c�"X���
Q�!eXz��y�;��<�VVː������T�5�woI�W��$��iM_��j���V����>���T�q�����������"��k$���)�ÏZ� �)�΀������u08Usx[�J�iQN�a���e�L{_,�o��sjꋩDD�M�>A���|�ͽ��$P�(��'�����d��	�BI/������e�[d�����~��G��7Zr�	sCk�`���\=c1Z��J~�_�xۆ{���6�$�k��= �[1ng3/�7,�j.G;[#"��2�Iy���	�ܝFJA,�t��֤C���\W�
�X ��u4,w�����vl�Z��86!����e��Rb<�`�p4���{tiN~W|��:v�{p�a�V���!c�Kck�UşD�_���
op��Q��Z��T��&��<��}������qQvߍ�0^^�W\�[K�����=���'���O�L���*tnf:�۔l�e$U�&Uڷ��V�v��-�����`ak�2�G�l�
��M#8�h�[���� ;$Q#h�o�����#<n�&ÀV�]1��xu�o@ED�qͷ��r��O��|�>k�N��y���nP��-���/3���r�N��s��qN��C9@� �Ӄ45��C���P쓳��Bȓ����p�'�h��&K���"xGJC����a;���H��Ѫ�+����
�2C�7��l$��EU�%��$��aqIJn�'�HsW�v���΁OY��*���ƍ��K�0�l��Fn�YOQ�.m��O0(�n���ϼ����nG���<����h�;%3w���3�}��8l�cJ/�����<����
�q26n�W�v�e�>�g]�*9ج�?�{�=��Δ��AM;q�-S���L�~���.5TPA�!��4w9��N�&`������ ��빤��S�`m��`�G
52��XZg�,��SK�Rl&����}�b�xy�7G�iv"o�^9�so��������&��R��d���b��>�9_���O�zf&f�&["KRh���)��k����	�uJ����P� V9� ��g�1��8��8fف�976�p7��x�&
��]T
�6��F���L�)xJy]䦊��)x��ry-ܷ�YM�ň�& .)�ګ�{�A%?���|e����DVj�u�D�F��Kf�	�e��O~����K�N�]_���d\�!kk% (���tn����`��ϥ��QI��9v��_�������s�u��5��Zc�AB"׾4Ciϔn���n9����o?�bU-��07�j|�X\e��dqY�k$�8O釻y�an^?��PB�0��8@\[͎>|?`�\�#��c{���%6�a���<L���f6>�"c���:���G�{��D��y��W��h�2TK�1[�G��a��Pzu�5Dx_g��M�i�t���ɀ5�'��۞TUP^��� �R�?���|p,̀��32o,f�v����'v%���g������J΀+%]9�+�[v��v���8y�F�r���#��?�朏tc��|1�Z���=�'A�Y�B�$z�xʚ�Z3�>ӱ�'��C���K�_\6Bs���<�B�I�9P�Ce���zUWgo�� �p!���հ1�̵B+o����4O�R��|�}�Y+w�H_.�o����9���5���s��k@S�h5�>ʀ��fԵGl�"`h���wlyN�QRM4��Co��R�1�d�}��Э�)H�IF�sU�y����S�MH{��~��h�d:�k�sX��[ �Z�:��+a=$r���B���dg��2�0���ՇB�n0r����0����:$���3�I�׭KckG��e��|>����t&��ч��-�I���z�K����[� ���S���t��SHM��"�U�C���v�I�Qv�U�;q	�ozi*i�mJ,��-��+;*.Xϵ�ɶT���$u��d�4@)A(/��Pqx�.(
מG�^.��@X@�?���ֽ��^�4X�u���JIv^���NA�oN!��b���ص�!�ĸ>�z 7�Y��:�ЕŤ��{S�1�R�w%���e�!��/�<�y�����X�;�,g���Ov/�$l�wf�����\�3�N��q{�6G��r'�l��D�oQ���owV��u,�DҞ��KrF .thW�Q��K,9�F���@L�#�;y�|��禉8冒�S~ɹ�x�r梀�o��߰!6cc]��t�)��<$�7���8J����M۠��>4��E�l ����pN���V9d-��&S��'�I�Q��T�}�r2�݅r��@���e���f/e�� H5��s�;%Ԯ<�(�������!��b#܁�@Z�*
��򎘊��#����O�c�L���y%oJ�����D��1��Ha��fMX�@�Nzȸ�a����	!F��¸PDe���i�+��i�P�dL�S%4s�ai^�g^�1O�����w�$n���jt��`�X��h��W�bp7N%�Y~Dƪ��p6���Dt-sO��,c�8�̯'���y=���S�V���Z�+ ICH5f��р��^�7�=�#p �L��U��6��~Ӑ(ޣ�*U:Q��7�!Xk�G$ ��h₴;jK����_"b���wX?4��%�D��5�p�\J^��TM�Zf(	;e`ͅ����p�?�V^wi!ԝ]@�^�w��9Ηz%��*x�ҖJbj��/24f��ώ_$�sA�JU��mx��'��&Ap'�sZF�Oj�{��V�CM�Y`b@�5ҳ�Y�Q"C<�{��5��:p��������yB��ٞH��F��o������`���q�c~M�2Lh��Z����0�b����3��q�#n|�r��ܰ��S�U�E���Cw��ydv-֡C�1Q?���ь4[i�}��R�ak�����9v}��x�_�!��π��R��DxF1�YϮ��/�g� ��:�v��]K���"�[��� ��+�\��a(�@D�MSbd��w�S��EY`#�_t�j���^�	�ys~9�ݫru��>�.�*��n
��|�G�ֳ���3�-����L�N�ߦmb���q���8�\u�����\2���9FƼ��� {gN����*fI��gC�����^��J�ף:���r�O�����ǁ��{��B�[ =h�GI���1��s=�߇�� ޭ�g�[����_��8 �2�k�(�*����y��tj���+ѿ,M��K��h��}�a
1�"�|��bٖ<�+�83.�NL�SR��p㬎���sY����a2��K��4�^�ۜ#�_C�"n�� �v��+^���6�%([ �i��_P�k��gU�t��Q++pr��z�+CNt(�Os���`wc�=p\��79`&�ceN�eC0܅��&�Va�e���GhdJ���lΟ�W&:�k8l�T�H�� �a=���uώd7�����xV��"Xi�B>�1�y�A$�g<*J����CW5v�y%X_�>2�5���(/<��d=(r;)*�A��n�V�E���p$�[������O^m;G8��*�/vc��>���|0��U�[�II��*�kãZg��%��
�$ټ
�6?K*P�_9��5��H��8��^1C�p��D�`�u�:��Ig��康��*�P��m�� b�,�U@%t���R�tn������̌����"�̘�a��*��0�����.21ݯ��
��P�]����^�I���4Dr7*��˦ e��h��r@0������+�Ϳ��sy�ys�o��\^�=��jHZ��в�	�qz������1�6>!�e�/VL��c��t+~w;7Mߥ�ko0��g��L���Vb�8����l�Q�
U�Gpw?{�Ө���j��\�%���w|�3k���"���$���bq9 b��h�S�Z*���t�T�/Xכ�'��ꄲV��Ӝ_�d��Ť ��X-|s�r�v}0�I�F(�פD��R���K�o:�t��L���U �8:n�`�8_H������1��g	t�X�0��b�t��LXD��Φ��1��{�GB�8q��0��H�yQ�šr���s��(�n
Lo��oz$�8k�PV�7�a��˪���W�d�O��EA�ɲt�~٢�꽻Y�!�o�#�l!:����(�RӀ�؁���!it����l�>��������;�Q��P;M��"6d�Q��n���F����Mz���o�2��R9eé���f�9��$4���\�o�e(�����,��\��g�[��Rs�ש�X�O1y=%#y1�G�8�L��_�}�I:��&;��n|��)�N�!~{"8��xe�d S�1��v�^Y����bixe� �30
dl�1���i�e�����������#cHF&T,D�m��g+���g͒ ����f*ʄm&#z����ܳ]�l�+�� �g*ªJ�cΖ}�o�������~�{�Y�S��&�����C���d�.�~��ORX�����y��L#�	�LW�$L����r�����rrnE񉏯jۖW���U�N-GTU�&cIk<��9Լ��\��>����-8 ,��fWV#�|O���8�<��[��{�x���i�`o�L�dH��ʬ���b�u�'7V0t�����E���G�F燠��o:��r=�˿�<�U�[�uz�(�f�5����^a��+��!ii���A��:!=�,�	����TJq���<!!��rq����yo��0WE�B+w�-�x�I�ծX�0�������w�|�e�AFR���|������N��ܥnۥA�ҡ�b����J�'�	���}�[-����٢t����ߎ�����Z�0ױ�K �f+\��ݿY��H���D"&���bG�=�`!��hǮ�	G.>A�c~�\��E����)�[S�;	��\���{+(c�D/���9����Y�YOA�_��CG������Q���A��TS";�t� -\+��8n��s��s4,�!9G�+>�v3��1�B	ʵ��]���,����ub��8d�[{D�M�֎w�F8	����{����d�^6���|��]T�� Z��yuIx�F�D	φ=��z�^�K��q2�SQ1bL=r�a�F��^m�
��<�e�	����m��C�@�Ht	������m��v�`V��P����њ��D�X�cwP��<�����-�ٞ1Dxq�;9�t|H��-�J�L�]�虦���I��V��4Yؗ#[��r�xH՜<.<����@�^�Qi-2yi y�t�(��c��\$zgHw�tCh?��{Eٙ,TV��_�0g�zhZ�u7R\c���-�G$^m�2�Cx��[k�<��L�n[����U�|�INS~��E�/��/R���ӨH��|x�u�ʷ�c�R��[}�R�v6������ޮ�q�"w�Bl�E�1/�I"?�.���~�W2xk[��7��k<6�}�T�w��]w�_�&��RU6�ܵ�Q���;j
����\F0�`�v��l�V�����ޑ�|/�8�3�$f�yҒ����W����Q�H�\�@T�ެ��E��t���{O�1E��Ҳ�O�pZ�9�0z��/�߻�!}P�*��ǘQ:��f���ei L[*ʗ���N�j|�p��XU�����m{isI��\���(��k�uO��]���A��9����dA2����0�5�j�vf��w��MG&n��b�5e.�{����o̯�������c����}�,���:Z�Yɗ^�'CaED�^��k����BKޑ�'���诛��F�,��[�@������)j�7�aU0!t[�9���^[�+�х9�ؚ���%>��A�t��⟎�s���s[�KQ�"�L�bR�0�K��J����s,յ�k,����酞-g����!IL���>#�Q�Vw��jڳ>���Hs��e�^��1%ܟ�+�>�!�	y���>Аz��!�!=�9�R��JR$D;���9�����Q���-i:a�؇&k~	��6�U�\�e���&S[F�X�wD�қ`m�0��y!`�]A�F>����~����v��Ï=�$�x��yS���/��Ǩ����?�����r	"Iv�8��*�H?Wт�^<���д�^ޙs��Z�#�'bR����n�(�߼�r	s�?<���5��hg�����(��$%Ub��\�L��8��u�S�PZ�!j�~�J��EFE��Y<��b�c��s�\B�K�A
��"���Z3�)�)]h�1��KF(�mhڌHq�.�)�3N�d�ot�����=L����4��Lr2|�jq�-J�Ζ�8/������IF�0�!Q�4��J�T��������L�
B�)�`H���ٿO���=iu-\X��+_r���.H%��uo<�6P8B�Lr��$S��O��>��=��s��L��nO�P�0��V]�x,����G�%f�u���5��H��as0��Da��a�{M��]�)�{z"6 ��8�<T�ɱӹg��Oo����@-��ΎE��S�~��2�Y�<(�J�p�b�D�vP�^A���jy���¯����}�.Z~�2�@����k�YP:��}A�9�_ܓ5K  �ݡ&�6E��}W���ehL@�)d�Ӭ�:Q�x��W^=� �
=ȶ�n����������9c2�������&	�P@�=:/SxT�)���cO���vF،�t�.�����e���8��<1Lp���D�x/�jV�~KY>b+2�6� �T�ml΀t)��`F|�oQ@i�]b���S�l���1�:L��*s)���aG���V� ,}����LLqS��&��}��`��)jb�V@��]�D^ V?�/��q�ΰj8� �ǐ5���k$�ߝ�m��|^k�m�<�p:��Br�Y��:�~���;�q��
�=׎�ϒ����meq��d�4�ʪqk?�3(\lc41�:��h�x)3��O:s����Q)��I�4�Q�{�W8Ͼkk�!}IJP�y�m*B�\ӭ�1�I��TXTFݞK��)G|1{�04�%ޛS��ui�}�F���#9�M��@�G�$P��H;���1]�]J��n��Nf�����6Q<�x&���:����]�+�v\�@�� A�!K�qM@V0Lkۘ}�>'�Ȁ���MĿ��U1oN�SV��x�s�Tb�ė$COl�MԴ���u f�r�ܹ�5
��lG��������
'���B7:�����J���M�{1O����|��Ln�� �5ܥ����n�WU -�_R���ҨV�C���O4=�Zp�a'��G]�,����R��X����s���	TȈ�I�ҶN@X�I�J�Z���ܝ�Ċ�F������O]_��/k%��>j,���F�i⍞	`��4#�1����.�νןǍ6@,�B*ٖ��5~(Z.(���uI�д?�.E�ߔ�$-��@��Q1!_�#v8(�w2�"��q*��aZ��ۍ���-�*��:mm���22W�T�#5j�:P;,��"�"�<�N���}�fPo媴`H��������`Vv�8	3�����;gx[�����惢��G9qb8
�X�B����������["XʴP�����Kt<p�ޠe�b���Xt�W=�a\&Q�	w�r�F�<��܇M+,a�����c�Hd:'0 � IY"M�qVFX��j���#K���ŗVQ�������u<f �x�#�[w�]l
�D�b	]A�E'Er����9|Ԩ�cXK*mg���pvy��)�>WoTa��2 &E]�v�iQ<�G�!�������6f�!�=�%����B�`e"�?1ԲN�'��/@�8W����{��tX�e��-n��6��E�A#��6��n�E�W����#`�!�*ǶR�3o��9Vʁ?Ɓ�(��٘J���^��%�lp�hw��sn)Y�X�X}\��p�t>��1k�a)$��@1�?V�^��[�g���M������ 唡a[y.�nШH��@�/�R�������'ڨk�T�լ3�Wׂh`��b`=\�pL��l��p�X����9ڑJ�����T�E`*�[(31�Gҭ�\3���A|�w/��ᓚ_�`woԒ�h���_2��7׉������]�K~a�0�G ���+߽x�A�O�c���v��L�5!	���L"��$W�	O1ttڂ��0�$ ����u�Z�0�l[/I��J��)r������08��.Lg_`?}�6���θ S| |��lvD���A<�
�Y�od�P����R�I,^�	ʀ�}c��BݴI�f��/���d�9�!m���� �R��oE�/���8�/��tZY@<o�1�6=��,,������u�S�x�O�Z
�N����ʾ�T�ƃ��T8Li�:o�ir!�	��3�1�g�X WT4��O�w*�_�#_ ���H{`K��Ĺ�'�|�'�R��<�-'���X9t���4/�Gۉh�e�z:φK�B���6C`z�cguXI��q�U <���6PzמUL���J!Ҵ�

�پ�%��'7t���!C����|NP:3'@tK7������DO/�l&*{7�=1I���p=!�G���wG*&�	Mo]��1�=CN�a��S��H�-aY����wy��8����>���_��k����Z&��e�=hP���	|  [^���k��P D��C�!�ܔ$�t�	���\Yi�r���yh|XfXF`�!�@ɀgWp��F4s�A�혘N�x��D��]�m���!%���dU`6޳n) ��!���Mq��~��0�Fy�� �;N��ۼ��m�ڰ�}RH�x�d�����:&B��O�|[��D8�vJ��@���I�/��g�*o�ך�7�̡��8+�PF0o`�e����b7��9��-؃QhA�)�n��{ĥ'��H�8��W��	����뿯�>!I�.W���[1��p�fY����;�D�
��z��-� �d�)'�m��I�\���-�3/!!���Wh��7��H��C�֮�vq��?s��Q����"I4�7A�2��B�OT��*p�tT�o#��NTf�z@X���eP�1t��2��+���'rw��V���3{z�&�e��ߕ��7�z�>�׾~��p��TCQ�:�$}8��"~�l҉*�*!��)��ڥS�އO�������!(<��t_�k�($����B� ��R���r���<(sq�9T�-���S��F��a�bi�z��M%d-M�׽rk�:�!�Y�xd�9��������\��y*|d�J���D��ؘ���^�gGRD�Z�#�5��,�����ZI��@������:Vl�J��9c��}�~����U�G�7��,O���^�7"|�^�$�č.��PnO7ɬ╠D��d+�w�$b��Ft煯��ծw�h��!��IY�ы�+\M�/�
�}'���Q�p�����Z�
�/�Lf����,��K k9�06���hܟ�xI4���b4X����e� :(ڰ�@=���1��|B?��g�|1��Sw�Kg��j �'�x�.��TKm����|"r��y+�u�3p)���8J�oH"U��Y�Mg�Qc�mS��k*�3e`xD�d�˟�� p\�_j2�<B��]:�=X�(�V2��g��@"���[�}&}�;��D-�-ۋ5/k��n�D;��HL�l��b@Q�V!4]�z�t���_����7����(�fL���oR�$�	��"�,~uxջ6��@J�-��G���r�Nu���eϵ,�U�y�%l����PY�O5:7i���U�����~x�mb���L2X|��&֭K��w:�ϛR�҉8#U���!y���:�g���#Ɏ�&��.�B���lꌏ#����5ԡ�M���:�/������B�<LT� �9�I����p��b��aA���^
��|���:���2��\x	Jtw�U����\[� �{-�mY��o~�V=����5"�U6I6&^�+?|\�%xsYm���F6�x������7����_�;��$�Ʀ/�5
��Xqf���O��[k��T;�H��M�Px�N��^d�USV6��1�,쳣��4��R�|��8i�&��5FSM
�g���</�wy����l� *{Y������^m�%RS�N��_��^��1�&��4�6���bt�s�6"�+�a���ޭ��j�Gt��[�jfKm����������Ը�3��`�jH:��I	*S�kǚ/�x�F�#*��Y|ՖG��Q��s+0��O�p�Մ��(��q�D�9���d|z�QL�I�'�Z(���O�aZi\P.�/%!.���3��駡�]e�b�21߈��L���O4x�eFqʫ�З����5��<�QXn/Q����O�tJ ;����p��		`��q��u?B<�/�~����o����Ug<<	޿o��|M�*h���Z
�Ӄ�9���� ����K�>H�C��9ӰUT���Ů߃���(Y�1X0=��.�������yy([��޽Gyf�Mp�ZP��$�7���t���y��=h��rxEiZ}���8������.a���5ڄ_��V��` k��D��Lh���
�ז��2�����n3=P��Y
W�R���1���Rt�zZ�p���!Z�7f��?
�%TVѦ����8f!d��ʟ��%B��+����w2��}�� �l2
'�d=� 2��Y^v�j�c+���튵[���������y�����l�	S����9�w�yZjw~��J0��vTw)����*A��˪'�C��͆.��)g�}���;d��_<dS�6��+��4b�D��4=f
P�x��A�����J3)."z3�܏Ji�]�ԝw��Dd\�R˟`�c¹@���(�@C�.8O�=	q�����[�?�͂�UIp�d��Tf�d�iۊ�֖�X�`�Q�Rم;��_���ƭ�Hv�4�i�jz�#�4�w���mJ�U����LF��"�`�q�R��_���	N���%zЎ�O�c�h�L9v]���|9ήd�zt�H�	��h����5J�"�*nW}���7��)f���y����b�1m�Τi���z:�����  B#�eWn��=B�V�",}$��vfO�㋃m�q��X�T�
1��qp!��a�dt؛}}\�V]���f����a\��;�8����t�}m,g��[s5l۟��h���������.��|@�̈�H^.eպ4�@����k�/��{%�j�˵߾�*��&��0ￏ���p��:?i�{΃���-�	i�����?�h�w����MCh�DPx�����2eL��N����-`��_�[����\�p[�lKn}�G���}��L��T��o���[;{EÎ|��ɳKFb�� �}�Y�F>����&�5��il��j�ʩ�e�ϑA���0�#=0�'�n�L�<��7"�!�^ޟ�K9�,�ˍ\~f'@O�v߷�g^�����-�2#�4xd��;���!k��R�ط�����S�9?�:���q�n���:��u�/�������0�����8i;��\Yg��	����q��_|Y���QϠ��Z���g4w���.�{�q]7�Y~%��C���K�s��}����7������(Q
JKWj �DK��V��CH{|BB��+c�W����#�t��⫣���?�o1i�u�B�Sy8��U�2��c�l�ڷ�)a� ��0�ZG-NP�<Qmy�=9���)�M/�zU��Vh����:�����.�#���.�/`��N}����k`��/���a���U=��D��AbbaG3t\�����;%��3�t�UF(�C�9�B)� �fL:MA���ho��Cx/����X d�}�������/PǙ���bU|{ ��2�'�����!ۆ�I&�Pٗ����Ol3f���]"����1��?{M��j���u����b$|!]�ff5�����lӨ�_��+u�.y��<����/c�9-��w	D��BT��pq\�S�uש�u�Y�	G�����]"���Mn~�-�D�p?�ʄ�r��+<8��\�+��4
�Z����"��*E�Q.n��w
���iF� I��Vo:��&�v=)�0Ip"g�I�����0z����_B�E����Y@�S���B�߰��
x�q�)W~�}1dY�@�{�E@�"Xܡ
�§� �c?+�ִ`��qR�\�v3����hb?Q�B�^2�(�bBlK 90l�7,|�x���/\H8��Ɏ��
(+��6��'��j�) �-݈��A��A�fP]��nl��w���מYC��������LU��k�[��uT{c<5@�H�N���<�N��9��y���I'0��E�a����)�×�3��}B׉js�bq���
�'�x�����[�ǽ%Q�g� ��r���{"x��zW��M6l�q㰎��S�.��{8TL/���GUWsZ8�Sh�������<���`0j�#_a��aT��F̼��}YA�� =��ĵ�#.�{4GSx�{��ghѩ�cY�[	���:��d�^��7�i�oq E0�3�R	����BM���ܗ�����E����&�����DX�ˍ�ͽb�V	_Cq��<���LsU@?h��g��7��U'G. i#:(]K�T� �g�@��L��q�S�BN�2,���&���'�J���-,�蓀YS�����!�7����&��v�ݟ���$Y8p(�����Z�0�'�yu���!?E���8�!��kJ�X���$-���4D8�;�r����ke�~>�p�T��=a�<Ж"0QQeA5�N�6�%�� �����1z>\�gw���y/�K��q�z�=1#ގ�^d83�2g��vG�F.C����t�{��k����_���J�g�q�3!�	%QtR��f�B�&>^�gf d�kА8������%�K���hqťf�*�q�Cb���F����{xy&a���P$Je�A8�����iGk(����y�,���o��ڷy����9�fAD8���ⷤZ�jꓲ�;)-*���y�u���w�Z-9ۦ�B���ne�����'\j��h�F���{d�֡�.��k�/)�A{�+��QE�y,����f�w�����G0(�5�m@'A��kL=e����t�+���3�3��r���̡π*L��s�c0�N5�ޚy��C8�s9�����-���,�]�1�C_���'�Q��cwǰ����N��<�1Ǿ��t�m�C��W`GM����KĒ�@��j	%Y������f���r�R�+6+���/0��,��[�r��ٳ���m_��8���J�s����M�&�1�$�4u��ǩ,�n�G����;�l��m����=��{x��ۦ��(�x�"��Y�~� ���=њ;`�����"$ �0*��B��Xؾ��FՄ���)u���*�^j�	R��e�������;Gp>�ٌK��Ԋ�j�G����,6�6d���^��Y�󠫎�����Pق�)�z�^�X3�9�E�J�o����-]��X�����hZ�u��k=g��#���j��g������|I&���P^i�J���m��|�v���Y�)�*��e�Zl�6Lb�c㦂"�x�!��I�pY�=;��\9oUV�C�����\$�~ �	鋐}C�P<=gS��![;�Z�����7g�\�>pP�_�<<o=��d�Om��|��aӳeڭ�뻴�����"����ͫw���S�$����(�A�������Ydk�U^]�Rة4��)��D��g��Yq=>zP�p��=;��U����?��S�վ�DHe�tD$��V�T0� 
v+���7�b����G��BxQH/A$풙%�Ϋ�,^^Ǡ l��!�C��UoH5�7$�ͪ�>U>߯�ݵ�d�e������k�l��@��'�_c�ƪ宑2fQg���G9�i�%r74�Ay�#�!�X�QxwVa���������MŘi.d�e ��-�{���-z�@o����v�_l���D�Z��p�!93�x
��
U xp�!�]+Ctږ��E�Yޓ�n �
5�*u�=�G9��b 堘��!�f����x3��,���M�#�a P0!o��jľ7�6Rr�u>�l���jZ�y�OkT��hQv�9���pp����ȧ�����#�Ə!1�Z�x0��fE���){��' �S���NĹx�����"Z�U;�7p�߼��F��]�dG�� �v�V�[(���!<(VB+��t�۳(_dz:�iP���<�\�!����F�4��pQ�?=�BP״Pw>��!�M�X��R䔹$�W��� s�!k(΅:I�w��^z�"�ʯGq�)���Bv��s&��⏙��֟�
���ְ��"%G��R����Au�z1Nru|&��!Z!��r%����A����(�r@q���ʵ/Z�pA�ˈ�ڏ{&� _'�z���D_$\��i��<��؎�"���b<�p�)C��4�����gl�DW�c�șD���p,?� �� �Zbz��a:+_R�
�"��ED��²�G���	پ���x�>}ٽY.9�'�:M��6�}��������܍�e '����{c9����&`r�Btr�a�X��4:���5(7��Wa돗��#,�%��J=�>b,�ίnI�c&���BO>���W��\�$�y� ے�	Er�2�\K�p^&����Ag����ǒ���_�?riQB�X�Vr�%��B.�a'gM�WV?N
�H��ȿ��C�ZVpl�~���p|���ܒm�۱A]|= I�YHr�*wS��u��(���[^#=Ә|�9f�gg	��e�e���6.e�;�k��'5|i{*���!.B���.�8)�sѾ8��j3��k��$c��@S� kŴ�{k �@�q���P3�Mf"��V6�Ob��!�k�LS�yUq������e����]�$>����(�|�]��$oa�S!�ϯp�6��.ᚺ�&�	~s#Å2�	&���+#cT=������k���' _#�#���AОJ�@̀���<!\؈<�)gWx_�,tS�1* 2�%ۧ1���Zk�s3 oH����"4��/�����C�$���ŗ�FPu��|�����_�m���5U�:Y��]�l�fzT��=�xպe��� .3�.�ϕM�LFL�|��-NԻ�V��J�=b�w8�x��������l��KSc��9	��Ώ���j`8�����=�6t���%k�c׆����>�u��O7��X\���͵%�����~u�v�|��p�-�L�f�`|�$GO�m�Su�D�c���e��i�Y�Ele;��<�Պ^�*g�>�d�t�&0�R�8f�����C����Z��6��QO��Tr�<�3�\O\�بuo��;���"L%I8$I��!��O�(1�>_[��F�G>�� �ϚI�Y�^Y�;#�����f�k���
0��lً�J�=�B:0���1�$�(�V�g��!���&�&QSc�=s?��1�}����.P��k��`�g���72�n�/>I��4�	M��"\}�{1*ᙞ�N��h��Ȧ��{,�����$o����p��c�d9_�K	.x��}e��`�^�S�y&㖫N̼�#JY!y��1\��!lQd#������B�YBD�>�נ0���Le	~�l��Zh��[H��GrW�/��?�$z
��֤dy7��J��#��z�9��{VW�ZX
u���4��{�YiL$v1�7CCGU7�O=�Z�P{�g����d�=��}�7�x������΍�Աm�
��8�׳���wU��Y`m���56Ql�$�E�Z�޶"��U����a�t��n�r%�S>�+R7q��Ո�/�	`�^����=�RH�@�j��.H��D�}Y�]3����d5�љ���gP�����s�sf���`'�'���>�9���c9;�^�B��)|��aWV�����y���i��vN�\��dG5�r���|��<��_S���������@��,���hCL���Q����@��m\S�c��:�|ÑK]x��C	��U*g�/=�R^��m�U%b�b�s���8¬o˿����V ��8��b~�W�k1Q �A�^4��c�^�,δ9lm�\�!f�\��?�'Z #��udُ_G��א��L�#�$���̩��FӘz�~���Pv|����ġ2 �w_i�����^\D�3� gg4�=9WJz�y�Au/��I!��4i�+&v�3O3@>��0T�(9�R}�獠�z�����$Gf"�Cr�G��,N�nEt���A/�|�cj��#���~�KQ��Q�i�S�&u������尳��!�6�kYg�
��7g!O7�(��X�/?�w����f&i��4��>�E/0�h���`�~B}���ʥ��t4�/�r
]�;ƺ{ujb�mq�W��� ����C!�f��W=�-�S����S���S�eg[��@�ȋ7y\�������ZK��H�e�����_,Fe'�`�%+��Ȟ|�V �mM�;��5|B�o��?pxJ�~p�s���{��A������v�9��l��b����mf�����B3����@�*��Nڂ�����֒ls3O�I({�Tg�,8MPj��(L��,�Q����>?��{$���D�,�vuwP�轧��� ��lю$��T��dY�Q�L �A��b���*_����#^`���	�(d	zvy��h�����<6���?m��xN��to���,����V"o�T$q��ZZ�t#{Z�]�\���r��+�AY�(=��<�c��G����۰~�֏���Z
�IJSFY����3�Y ��"����{�-+��6}����Bڲ�2�^��n6{*����:od�����]u#��+d��?��M޲�c��-|)Z��U�~�
j�^�Z3͎3/�}��u�}�a��Ǳws��*�������[
�</x�Xa_�3��퓁��#������Č.�N9�������1#H����-l�O�k{c�U����e|`��
!y�x!����R��t��I,n=�Td�d6�P��V�.8���[�0����?��o=��m�����U  a;��fԪ�����2��7L�Z��3:RF�Y�&8|����ߌF�]��=;�f.[��oG����q�U��|��蘋��&�qR��<�l¸j!X�)[*�8gK�Nv��NE����~m�~���6#9�xKR|�E��:H��e��K�BB��Y#��*g���DH^�-�U�#���.4}��n57 �@��x2!�"W<��a����g���?a.2h�w��Ƣ�y�7���s�V�#��Yq�2�+��T�BЄ�n('5�RX�_fo7�'���7A�el��Mm��e���eٮ5�aK���N��[�]�
v�j��Y��3f`��h���9I�����e�X�YAg�[�4��-��7NBN�mX�b�:�+����ӛ`O���Mv/�eQ8�A����/���z%O0^AL	=��R��%�W�n��9/�91�-�+�#%��%b��ܯ������N]��������/�ݡ�F^*fͯ�p3Y^��DF�y�X���fj��1�37�W" �5n��¹M^��I�|w��0����*d���> ��R��R��� saz7�j���.�9�L'�?o�
�3<P>���+�q ���}�h���N��B�(�*%�ۜ�4���gy��_m�&u��-��,�~���u����*W��&��t�����w��A�	lƕs�`;g%�yp��������P���o{�ok\ϙ!��:u��S/�F�[x��B��ק�e���X�;�cRiz����w�Y���x�W�ji{����!1��M����+�N�h,6J-�d<wzc��i-���@o�bx`Y[�|�D�Nh�\"�?R��C)&[���"�hj�%�~�7����iP��JE��GcW�GsT@T����5Z�C�0�m�f�����/Kю߅;���������?�{��Q:-�E�ib��"�mg��#k�7�MPϟ��J��&���մ��%=3f,L��Q"���r͗��E���}�%W��Z���Hdl�A?�`Gߋ�����&��̉�k�K�G��Q@3�����?zd�@��115)� w�B��K���ZU���/��:����
����k��Հ���1ȋ_˙���C�p��@��R!9D��"E>���Rh�45r���	ѝ��$���S�Vc�"Cӧ�[?�L�����x��E#�et��ꭓ#v[P򊏨�:���<lN"��:�+IMys��m�;�TZ���}N(t�޺<�y�%J0B�Y���Vy}Zn�n�F�f��c�C���2!p4c��-0��k- �y'a9��|�� �Ė)B��e��o-�fʄ��n-ܻe����`Y2��m_ɲǋf��x���)7Qk¥�k�ܵis9�1����MA�6DK!>��h��b��A�~��]]>3��/�9+6�m��V��-����kIgxs�V�S_�=�O�O�b(�\��"V�I(+���r��9_�"��W#�F��UK�(b�Ӹ����⊡{�#��%$Ih'ze�-I��y��5og>� h�^��3�1����ׄ�:m�)�1���Д�ɖ����J���λ����-��}�9�����wC���e�f�
yoB��l(h��B�l�}}��j0Xέ�Q�V�>��oZ��a&�냍�6ab�w�
��Os�dxhm変1�Ʒ��ںb��/���]�U���Rh���Q��V�*}���4����;,2�CD|�mp����d�:�ڰ�녠F��$ʩ�F�5I������~l���_^IГ0� Zt~���1�7��:߆J +Cپ��.,R���Vؕ�DvyĈ�9��	�7��Lorh?w�Xi�q��iPҟ�y��X� `�lR����dv���$�,i h�p�9g�s��%����-���.��~$M����f}~�&Y~f�~"�\֍�X"���+��ht�Ōf��A�vW�bDuvd����SL~�W�%+��`͆7���ty?�G9���ĥw@B�\����9�'�rtw�ƛ�	�,9��^po����3w8���j�1�0iZx�Qi�Y�t�a���UT pm{�D�u�Sx2.�vA̠��0v#�uMN �Wc�g�(��&�QiӔ �L4��tW]"��|Hg!��-���b<�g����E6�m=���9j}��Vߩ(����#��D������n����+��ys#,z5��i���&�Z 9jI�}���q�b�A�K���x�|S�tQU��;��@��\��A~�>��}&�=���?2C)Ia�p�h	D+D��9~]��߾i�d	cUcvؽ���M�Qn��_�VH4x�)ڴ�[��-˿)Du�e)��7M��|L�Rn�j�h��9��I��Q�?W����&��T�j��P5�T�b�2x�;�-��x:�=�D�;(��U��߅��w�/�m=�t��ڙ +�Z�qN�7P��B:d���s��)b\:wj&�����pye6xr~A�hz���{d�LDE��م���m�1G���2{�{4�u��YM��KK���S�G���x������ ���1���@��v,���
B�4�c��Y�q!�,�*I^� D�h�~�(���1����[�]��O��<`�����Mo_v���MH��Tu���u9佀:Ɛivސ6���"�����3��\��;��.��-�6�RT��6��V��>ݙ8~�I�K�Ћ�	��L2>Y����)��+tr�}�6�(=vv>��=YL�!U�Ҁo��/z5�o[zmH#����HD�57'�>-6rCv���7��Kͩ�z���H)��r�Q"�5/�
�|9O�m��;�g�mHZU�H*s���L���"�9�2�'W��`O�8c�[�ScUe*`ki�?m&1r
�{�&qS��>J��"�t-�v�>\4GA� �藽��f�]�EL��(��e���K�]�I (by�z����F��ULr:v='µ��TK��b�:VS�[guAG�us4��1���o:T�+b̚�4�YҤ�{o�ɓ��}��*���Q�$�gG����mj<[AO)"袵��f�Ï���K,��s�Q��f�h���mC�d��g�.����s}����s��JdrY�T�%?!�hh�4ߙ�`�� ���;
�c�`�F7�x<�|KZ�i":�.�ΊLQe�,/��"�-�In���*�%�H�Kp���h�9���c}�0f����:�;�\nf���f9B)2�*�mr��b?�,�J?'�o�����)�(�$@Z���!�y��e.�������87��T��-����x�����J�� s@R6����c�~g?l�;L-�Hkq��}A��"+q6:�v�!��#X٨�l�C���L��V��3�h��ġ�W@8n�Q�(�P+9�Jo�螨k颦\ۈ��R����� �Ǚ��e�=�u#�+���a�= E`�e�ɖ��N㠳���7�I�v��ȒQX� ?�*Ƶ4���,5"�Ԡ��*r�z|��j�)���TĔ@�+�\�D�U~r�N�6�@�~FTA�X��Q��Ky�s)�����8�Dȳd��)����7��@�5�D�1L���3�E)jQ�W��2_3�
#~2١7C�Mm�]�ԔN�^�U��;�-���+������y�~�9��$�2g6�Ěϭ�U�A��5���K��du��#,�>y�︓N@���	�,�&�'=6��E�����xd�
�^H${���!�"{������������ť^���D��7m���il�ܗSN�<�sƠV�b��+��lJ�"y�ld�һE�7B<)�T�8F0T�,c&�CH�<��Ċq���7��C�$mɑ��J��#.����"���m�B�p�W�8#�yK%Rh��nC�|���R2�[haB������䴏�⪰��|.�5	iVW^�澞N�<�6��m��t�f��=��d�
}Wy���{i�@<��ǅ��!��|�>�QG�yy'앪Zt��B��/�i[�yY��mi�^"s�KF��t�R�e�2d�w��ib�9h�;����H��dn۩9<l
Z��Aö��f�'U�s�h������
���]E��3Y��ݨׯ�ya��u���K�.�=I��pX�ݴ'�C�3�b|5�+ ��V�����N�XB"�R:J_��[�Q�NC3�0;��,���s�E@���Z�`�O.���o�Xr��K]���;O�"�s�����^Lj&�.�\SaO�� ��zK�%)��F���!8�6���:��eͨ�'�DM�k�#��h�v@�*�?�5nMQKZ�Ӿ�@+=_Aa.˨�x	-�k�Ι��{�}�D���HT�e#!JQ����<�ɿc������{�L�ǛA'��Ӿ�M4��L��d�5H�H�8b����d��*�<_9d����꽎(]�b��2��A3�n��]��&�ʴ9���3�Ҡm��4�Ol����&^:d�>�۪��et����Z�kXy����A��I��,˘ҏ��l�+��ǆ��a4���>�I7�����mX��=wC `)t����.�ORO�/�6t�`9�K\�c9��3���ǉxVa�M�,DO�=���?#���$C��!Р���sm-s�$�`h�_1������T�j5��uv���5�5T�w􁦙�XR4��c�`��L8fc�2P�[M�/�(D|���Nqέ����ۑ��+�PVE�P�;��%}��ћ(��{�����Զ��ML��n����A�YӨ U�ރ�����r�ŵ�-�IOS�M^�#�
���בU���(Y#���W&�Xidvg��U�Df���pP�n��%�T���?C1i���"H�� ���I[
 �Ѧ�Ď���=�@���Q��X�Ji\-���Q\�a��g;Ga��.�Q��=�m����ZD�Ӈkw�#�"
P���6A���r�.�$�����4�����+�㶞kRT�Һ�<��i���v�(��%dΗ�u�l��o����,5���hx�#��!���>dh7�p2�R�]t�L0�����}C���S��Ց�
�z���Dՙ�=��o�]�����Z�J���}W��ɚy�MK�6�G�l��'GPY������w�L��}_��Q�!�0f��e����d�^(�_��+��5��q_?a����Ϊ߳Ԝ@ğw-��M4W̙���2o���!��	�W�
HH]!���S@����3�8�	6[�	����;�&����aq����k�7�[����	Z� D�Q��08Uy�A�TeP@����ᥑ�	c�qn��1\�Ӣo�83n��l���[��P�i����u��rr�ExY!�C�c�HF�m�*�U��pSxQL`�qŊ`R�wq�f"�;#S�� �RQ�sRc|-�n�� �rH�E�}v_� ���1H���5?n��77��T���G�-W�)�kr	�H�TEz�팾�ݡ�k�c����	k�A��(�ޔ�M�8��/=^�z���QOW�tFW�j��0�>��oh���n�-��(��'A���"�(e�&Wf�4탥f���������@w��(�P+	K:�K�i�wP���:爄*�2��_���,��:W��\�"�#�ާj�-Xz�1 ��$I�<!�$ܗK{���w�un4]�h/)����F��%����S6��n��HN�y`�8�6w�"7��G�G_�6�JO����W#�a՞��p��̬����q����Φɜ�.Aώq��!�+Qh��DN@Z���}�p�)�����8�=��D��\6�n9+��@��Tu�:}d-2�3�P���$�~��W�b�ʵ�'��ݩ�������p�>�Ƿ� ap�橙,�0+��h���H���ӭrfPY�Q��9xwM|0���8% �ʃ_�	TL@�2������,`P�r!��G7R�qT3/�������W�7�[�,S}� ъ|�a��P>Qy_��cl���8�Y��M��O�_�m���x���'C����'�����b�\���qĎ�� %1S���\����~����ص����f1��d:����	 �u�6�X6�D����n߫�W�aCH��]��|��t��p�&�O��d��� ���o�!�x������t�DO[�JS=�r��G��G���ů��݋�ES^�E�|�����6��k�G��FQgy��wN��A���-������:;d�l�F��3*K���d1���4w߰��Z� _*��߭�3k��u�ڂy�c"��i�/*��1n��,�T%�ۿ���!�]�'�����kf��-��ٞ#r ;�-B��E3BW�N������]"�BP��`�ܐv�)cg'7�6����N:-�	kvAx�ь���y�c���N*���z���
��W�u�W�	��<N#�<�M�����Ψ��(\�:���B# ϊ�v�t%�-[�U�C����j:�X.u�}�#W��Ri��;0�r97C�����㤴��
��T�-��iG3����i���f����␢(�</W���������YYSqƧ�"��#fB��G��T'FIq����-��I&%����>�%�MG�[�+h��ؔ��y�6eƭC����g'� �I��'��i�0��l���jQ��hE�]��4p亽�
95�����mY���*�߿����ue� uZ��g{��
��S^v��	&c�8:�t�@���30��wfW՚
 =8���ۍ�K�b t��%ԯ�� �L�p��	n@c��� z��Ɇ˄���
ۮ��Y.��9ܩ�H;����(�ʴ�Gg��cj�C��؁����$4�xT�Y�0����\1w��]N�b8���^�@y�WH�{� \א+�X�?s�K�@쀢�������Ъ�9��]:(
ͩ>$p�F+Uk��
vs(i(��D����+��2̇i��B��z3Lh罏�.�_�ߧw~���2;Yi���>�zfr5r�?q�6�S�˩�,���&�����|Q���@��N�#�$ѱaV���dq�����4�-Z�:{��fi�m���ڰ8���վM;9w	��S�i�����Jy#A��q�B���������m��Q����ѱ���5��O��#���v]��$�i�}wh�;Eq�/���4� �s������^ja��?�`\���Tޞ�ٓ�h-.��i��V��G�>�S	�b��}�L�&0'!	fe���i�|����'�#P����&�g��H���� 	V�	MQ;���JfŇ�m��B3��WH��Yؑ�$%|�ݻ]�rhɳ��-LC��D��L¤(�%�1\�$�̈C���
�i����s��3��G;F|���N�^�=�8��~@����[����ǻ���	���ㅡ�?�Ŏs'Qy�\y�����S�����@�o����U�����&#���U�����K�,�jf������9�u�cQ��R��u�&��`�<:\�oh�2-�^�����'⫧�/?�����Gvq���z�J�|�����^�!�vC�s��WC�}��S�X�j1,���n_��;�f0]NFMh�x����*b������D�N4r�-�Co�yi=�wA����X:���SO������~�j��5k��}��-1�r�����6�G���+ڞ�C� l�5��z��jnU��^��k���V�"�
���k�=�ѳO$y�-WBb!�	������b�r��h�L^��d[�<��܄y�Z�Ԏ.;��X�tj��X[k�pOQ���
"�
�՜�˫�������C���������h�.��q����M^8�����sUN�H�uM
��Ps����;:�Z1�V|<�c]+<x��>:%�dihf��}.S��ՠ��E2�W�sZ��`�9�R�����]�L�q6f�c>v�e����	���gy��:B`�Û�����#����;�wxc_헱�bѦI����^3��H�h̡�< :�_�H`��)�����p���?
�2�6�פ�L�nYZ�������YQ�J���)T|��K��NNZl�;N�֣�����k��P���a� �]	�8�jHq��S��$�o��.�_#^0��܎m�V�ܫ4#�=��j�.�]��v�v��eĝ@/�@��z�P���������;�޹��1�ԉ'E��'�i����W�Q	�8&�7�V����턳��#�r�~���]�4Z�T$�������g��g86��jM����Co*D���G���E����}?�w�9	�K��,�]� /�/�oص�u��A���nm;�m^�~�o��SY�fi�����Ꮌ��x�&uDg�$�w����$b
xA�t�c��1�NC�j�/Ojz�Z��uގ^�:���#�?d���0�$�weHz2�%M������Q��wB\_�_���J�����|��|蠑�`��<<�?��؈�q�0�����ͱૐ�s-z_6n�	�����R��wꘋ<rB�U�m���~���r'�2�L�#��~�g}�V���rš͊p{8ml���)��󥆎�ZݜV��:F�{uP`0�q���@��]�\	\o�5�቎K0������Gp�m'1���b�[��H#4��Lq~Q�h3$�ˮrM�C��f�(K������a������;oA�o�>9E����k��;@�\>_W&�1�C������)�R�����me�OMa�<H���f|�c�F�>/{NHG�nɺ ��+�ye�5C/g3���O�k+���=�� '��q����M��!�pό�~L����N�W�p �ɍ�ő�<�n��� ���>W��f{b�p�q�z�ՠ�6�**�-7�\T,�݄�w{	���ֵ~dLv�M������zm�v[��n.7U�='*�=��^�Sw c�ž��#!%xJ��T���q]3�B�r�T_P�0:�!�] ���7���cCY"ׇ�t�$2۪�n���j��X�J᱘v�(��T�`�?���f�\����v��4o�r7�?�r��y~��Hn�^t�>`�L~�I<Oz���GM7^�'ڥ�Z�9<ڱI����';��w���bT�C���C5[��1�ahv_2~�2F�`^;�ܻE�\{ ��H��:ȣ��>C��|�Q�an�P'VPy<�?�\���Fx��.m`B���G	���ssm����qUp����|�D�LI���UY�^�	`�]���$��2�|Q
�����W����Xh�gN����	��ge�(�H�ܝ�Q��gܞ�N;D�]դ�k3x����s_N���y��T���G�
�4�H{uL��$^�9��3��SHX��$��FK��^�(C�=x��zR�܉.@c�e�d7>��z����l�����c��%d�A�V�`yQ��oi�o1�	˫��Ut���x
�},{���amgEO6�m��гJa���i�V��(��G��=��>���?��3皎���@���K�yi���a����!Y���X�|�I)h|�$<T�Q��mݙ���BgW8�iQ�(#� �!0q�%{��K`ѯL�q��\hA���t�R��j��C� �dEĢQ&q+��?�,n/';5�r�օท�R�t�N�_�!6^k�`�rN��VUlF��1�23'8��oՂTZ��7�E���~uj�0�}؇�jx|0�����}Q;E����I�M{�!�;��k!��W��&T~��8��L�:r(u��i�n���w��.5����f�/��T�嬵����*���Y߯���Mv����[�xèF�bǂ�I��Rkf)�
�y��tiq�[ �i;�u8ҵBj�n��,W�\��w���tJ󓇕�!H6�� ;n%oס��ͨ�V����G���ۀ�f"!�X Y�d O1�")�l����~N��#WU9Z����e�z Xm@rJI'��u�T�E��:����Лa��'o�l�@��c�
���d/�O�*T��Ή�q'ؚ~���{�|��C7��0&������H�TD��k���+��hͩ^ñ��Z�L��e�:?���1�L&�h$R;Z���0
.=
z�Ʃ��x�h��w���̧�Θ���+�n�-<��8$��`ldU�3���[(�]��4�F�����,[�L�Xͧw
�'K���՘ˬ:���a�����$��>;P�/�/LS�� ��4f�rr�ۃX/�`EU�2!���PWC�;0}��Z�y 绨�#dz4�My���E�|FZcì��,{�̙#��
`�����B&	�������$�a{�g�0��x��*u�����-���?}���sm�(��-��+� p��Q��}ٞ�Y['hx�=�U5q�6ܶLR�ra�T$�uy..i)�xZVG�����8m�_����G�S��`W�n{p �c�/�������cT�+�!TR>�� G*'�B��&y�}�8��L(
�ɜ�J�J,��&�ӓ�+V������1��&�kB���"hb����T_x!�@��۝�+�d�W��%y��>�A��� J+<
Ae���d��&��*�����h����Z#4�+WN4 ��h���m2��p���iu�49|��$�x��c0�	J�D.���þ&������~�����>x��/u�D�@n�d�<��c�}�˴ӏ,��;4:IX���Ưs�s��hs��j��@��Ļ듴�e�׈4�*�bQ��{���3l�o�A�!0O�oa���Q&�ϕ�BĩAZ,��}�mr���J�q�{u��d����ej7��_�[R���t��J�	G����p���`�6��:�����pb�k���Q���{�Tb��������t@�B�A��{�RQ��v�/ZT�4��0,�S5�j����L*0N@Yw���mc��]l�{���I0A:~?���1�4�4L�"E���q��|�[R F�m��8麫=D� ��� `�����[��?i4�++��?�񳻄7�!�����J�ܗ�/��	\�<ʒr�F>���L�8k���΍�p�˚j���RwC��FrSm�C	<8�� �t�4��{�5b�
�4
9$�^UJb���0R�;��Z���'I_!�KH
����z�V{K���W"M���ZΛy�U'��t
R��J��Ņ�f{#TFV01�3R�>�zg&��]|���{h?i>%�hiM�ᄙ��&�W!bc��,|�8]�_-]F��5��#!m�z�e[���q7?�����s�C�R,�y�W�%$�[�z�q�\�)����C^f+P6�>>�-n�� 6=ʎu�PI{�S���$��60�f'�*z]��[����={��5����
�:{=Š��0��.�������C2YRfa�
�|����t���7 �Q?{�:k�+�D
W�D�G����z�c1�}���BY ���6��4��A/d(3��/�e�ƀ=װ�`�r-���xq7tV B�V�a�f�#�k���F�waR�n�����]��N;������#̣U��=;-E�2�m�����]��Qa1[��A`��-�6
6����*d�s�؀�4{.:�L)+w�w���Ș����@p�qSƾ���;<��E�#�1�^ނ8��O���QSF.��/v�yw��x�M#5OhF|���q�-;kV�����q�ꓵ�ui�t>
kG�ܒ��C0��xp�
#J�Ze�6
x�-A�)Y��V�4'R�|�eK�M��@	)��F�1��R��o,sPi��զ[H����y��_�y\�}W��P�	��%�mt[�@�;��4�a��`C��[�;�ƞ��#!�i��J�����)z:����ch�����q_��CcQurB��@�$]όGv�<>b�}���mu�X���v��+�D�����%O(�i2�ץ���$����f#��c�n[SѤ}�P�p�\x��[V;��ЭkY���٣��@+��T����E��u�p��0�ϡ�}BE��^ )̂Eh�*;�\Wv��|O�e=1��`�Ŋ���z�L�w=�vq�u� �� ���+���y��k<�;���w��b0<����0 $�@|�WOa����{o�ij^5�~�pG>fd��毝��ܪb?�;W#�0~�47����RmX�/�vNdO^i�C�����I��:9B59L"0�u��r�5R���߃Z���^|���G^?a~���$̸T_V�^|�9�G|{�<������	��IFxa���_G>�gj�;*�ާ�����P���^��)���(��Ç��5X)�%6��-�/W%,zi2����ڞv;�[j��U�7�NX��l�� ��F�skq$nT|#g\�H��P�/�Sq�{H���`��´��5rM�z(������ LZ��7�tQ����#|�a���dC(�����Q(�6+�܁����5� U�Ň�<�V����U��޾Q��S�A�������1��з��0���c��9CLY��y���c�;9z��~��({�m+͇��a|@$N�+��ZG�q`���1IҤ>j��^(��^�،=��X��A�̉/���S�&+����v'E��4��	�VQ/��s{C ��<%r�#6��3��)2e=FՑ�hd�,y��]e]�}o�5��燗u���ʹ���s�{;/��b�:�_��nQ�w�3������&�1��m�����ޝ����p���u#��-19A�E������O)��.ql�����.��To��͂׭���}�C����HsAaI�u�y�)�/P�9K���]��@���6�����@���`R5�8U�v@��B��D����_:�@Ç�{~�i$��Ðj��ïA�Ye&���aR���LK7�OU�����j�]��S�͜����{�gM��_��o��o��Iz���-bF �s,��(�\��Q�{�&� ��Ȉ���E�/�.��	]nnj���n�/�O��2ӓʙ�=��5����8ܛtx-c����@��1�+���>�� �7^�U?�����ԑk>5�嶇�D��H�^�am�Ϊh�=�XCw��D%��׮~UPH��^�ᝑkd�\���ێ�<�v8%�|�At �������]�y���~lmb��;�l��������;�$��ݲ���=8�Ћ�h��g�HY 3���ڞj}/;�W��ږ�T-7-ً�HJȶz���&�f�C\�#��@9�1D z����؏�<���[>�/�)B�P��;�E��)?i�)[^^�J� \����[�A8��F'�e��w\u�K��EʦS��fծ�e��F�&�k�XK-��W�C#[��A��.�1\Fd!
o
¢�ُ��\_u���bR��づ[�"�e!�����W�s����u�K����R�~�<}��w�cbC'�{���"w'�#������$v{��U>5;�k��9k�엁���[���c{$���R�o)x!Cq��͎�^YNlb!��֣���S��j7Fߏ��[DRk�|�/mV�2i~�anKz��8w��ڛ�����$�?O�}�xκ-e�%��Q"�`��G0���.���N��ͥ��!Fv
�<.ţ�ԲC�~��+��X�ľ�y�"I�y���VJ�/O�b�tS��Wevu�c|�JzG�͂ �T�%�묦E� ��.� ���2�.K!����~�v�~}h����}�$Gxާ��X/�;ث��vߝ�S��y�xYZƕ��9U�Cd,Q���M��_�P��ɿ��'��~)����߻��#�������[摳G�%�E�<������8ٴYZ�X�/�4��oyN�tg/�N����5�c]	���� 'Rٛ!�]-f�-����M)�Jԧ��S�(OT��)����鍐�J�Wb��M�Ӣ�h�v�����ii���t�O�f���}h�0�A��N:@�~G�n�Ny��"IK�^a��P&a{� 	5��Y�p����`��pP
Q`&�p�rG�NZ��m=_Ǵ��0���F<��|���$<]eң湵�,�I��7�P�Q?ٟFԙ<�غ�Ͽ���2 �}��]�1^��'wj�ֺ���:K �0�es����:�|�PB,4Ҋ�����������S�c����Ć���}�"�JW��h����1�&���^0��)�e��v����7_d]u�Z\�}������zZ�e��}[a��J�����O�H�����8�?g9?��J��u����@�y��,�[W__�Áy�IU-��qo� i����ȈV������6o�
�w�Hk.����1[A��@UYwxK���_�:/��7��^�ʎ�I1ق�!JD@�ܟ�H��}���%������'C\U�.#�ώ x"�0���L �6�(�`��G�>���J�`5�����[��x�����`R��j�eS�sْIO'�*�ve.FOD_'u��e��]	ـ�joky���/�m�mJ��^�k:�#Z��&4}��L�t�s4�<g�/�~)���-�PkO[WC��	����
(�g��y⹐�:���C�B��z/b�*�'�?����Ά�\������>�*����3�^�I�g˫�I>��H���B ��|���e��-�S���ZS[c!����&/���+�~C
o��b+� ��/T�	�����:&�9�������ϪV�T��[���!�Y73h'��%|��SB{�@W�� G1�N^�5b�!�<
ҕ�`���`�G؝2���ǯ��:�q��%@�J�x������9#��-��+�7&"��x�.)��]0��U~��9�e�UR���ӳ�P&Q������
�����Wr����jOm\�C+d.�e����ma�i��[-�$
��K���U�8ƞ��	^�LT�x��x��R>cϬ�����%l�O����Ԉ0)yɍsZ��i��|�I4ە�j�_�k�I�Zo���+)�`U� ��/8�a�����b�?v/ܲ&k~	0�~��A�3�o�m�CY�����:ěDz;�k۽��@p�%!�l0�z�:�$e�J������h��FP���|�Sz�nXT7Ud�!"7�R�z:�ė=Ȁ���W�b�D��0oc�r^��A�sE��qYP�\x��Y/�rV�Y��B����U���Z�}��ȱ�[\�"��S�^1HVҔ�����7��g�8�ڝ�R��͐�xl@�iơd��-A�u����B�����kɡs��c|j.��=V�W��G��Ҋ;��DP"�|��}�K��ԨC�F�>��H+�Y!�˩�(@�m�^{���"���&��i��΅C�$�~.�#86D��=�I�����3j(���КO�3;��-�&��EY��Ԗ�[�������6�K#^I�J
�y���#�<SQrJ�u0/�7��K!m�A��B�r[gX�����&_�y��psϚ�rW�^����^!=Q��*}�8:��mA����'����É���\�%ܿ���Y��c�������b%��H�ڵ�^G��7��߻�[�i�c�c3���$kZ�g�Y�9<q�^����|�!���l�2O��5�K�Hk)�`>r���gHI���)Wi�F���uB|G~����- @4u6 �?�&E������g@�F�a����s$z�h�!U�Tp3?+g�D�I)���a�֚�	yv���#Jh]}%��}�6��3��fI�'e�2�o��&�5*=�9�O��@�4*���uLtI�|�F�[U���R�|�f��.���k�6����M9m�-��r���zW�	�b���w�+s1㵯�h܂a��}�
fLǮ���.a�<cG:�4���~Е�q�<f9�m=;���b:�]MG����^t\��Hۖ��e����;��ܲ�=	զɘrG��I,e��c�3VX�Gj&&��C���K{��Q ���1u2Sz��`�B_�G�`=��n�܇��I����!;Og %�/��g_8G:�L�
�M��|���|����D0����I����|���K�^0Y��*��r -�C6!�^�hSA��) .Y���T��[��}�l4E�����Ң�Qd��UmR^�%2V.o�����:����[��>�`5�S���OJ ��<����T\��aIҶl�I��Ox���{%*��V|��b�D !\
m'b�~Veѕ����f����(��ڱOm'�M���H��[��
��nH�&��u�87�Ւ�U��SY��z�f�$깑��b-�}pG.G��J�W���r�=*C�4�`m�``i��Fn��ZiE=V�i5���ua���kp"����\<�����;+�5�;5��`O���4/u��wĤ��*��D\�����t��1��\�`$:9T�} �Y^��p	�T&&��_����������=�雚�^\������"�7�Qe>��n��Ґ![��N��n�½���ZlZ�d�ʍhRm���hMw�b�"E�)yk���ɻ Sp8��{�G��<,Ŧ���!�R�@m%n��>�^���t�8"U����W��E��@o����J�U�p�e��6��9���<����W��q:��[�ц�	bs�*7��(�V��Z��4���9�}a}�nX�%h����&�����9�ɖ��IN8U�؛���g�`����F}<�ia��|��*Ua4s�N�È��~B߾J�� �����(� .{��<�c��b�w\vkR~�SȜMC�;�o��^
Ex�#f�"
-)ό��"���7��j�W�qi��P��^D����P�����؈J���/1���!Z�?�W�I������o�{~e����u�NU�%�bk��3�I>*V�|<ݟ�98m���ì7�\�]�v1���W4#��0�}�Ȟ���=U�
.�~
|xG��E�񊊯��{1��Q�x�L�eAr}k��f�ܑ����_P�l.2��r�w5���Y�cv�u8`��l�,5�d��D̊�W��Wa�-}��>�K>Nv�8��a߷ڿ�Ǖ��ռ�����g��y�?���S�u�7<��bB���&�:�H����ғ�;��"j�1���+���s�co�F��0���'����8���l7>XUy��I�~�QOb�#T�]�B����)\!~�?��X3 kXB���Q�^�>�
H�4f݀�B��s��/���H�=9'��Ů��P�������/���}�e�^��p�/%�xWKe_!�R���Fw{�3�'�Prku_9�uJ�fTb9#H�A�E8@w����~t=���(�`�+��Y�����y@����+�b���I�|���6�|Ą?Z���g��9?�d�g��'��&���@�&��LR�1E�����#s��Ey269P��x�������Y03����t�,v��Y�Н��x�^mYK�n�2��kĔ��#A$v�lt��@�^��.O:-/����a?�:�y�����Z�*d��5ǹ@y9h��n��˽���+�Vz`�����и�k�Io�R��0"P�Nl\�Oa
���3�(�������{1'��=Nk��u�E�����{ۺ~�gk�du��`��<
�/���A��I�a�~�Y��#�D@���������Ի3��B?*y���1呏�>�(Ͷ�V�=���T��wmL�Ϩ�$Yl�>S��JLk�G�Z�Ŕ�~�s����M�y�~Fj<k��o_9�M=H̳H��t}� �MB1���\c����|���i�k��^�ъ/6}�uaU��;!kKlqf�W�y�}	Ni��(͖n2q'gf!�����h�������~�mG����j����I�dE��rz0�'Y�WBF�I����F�Ik��Z�~�)��1��w| �ﭧ0)�����m��[l�T"P��Yh�)S���m�y:$�J/ʭ�ԡf�1 [�ӴX���NT�X�Z�l�5Y�&�2�P^K����Ė��7|�a�'�����@x�i����?�V�{X� ���PהC�
��6�0�{<�x�gp�^�s��%�u��+n�H�շOY�������{��`z<��r��U���(�!D�LnN����0P"�D.����4ǩQ<ʶ`�v����b��'����/�ɻ����:�"����_��������c��)�U����د>�p ��	����~11���8�v��褈��X�=�0�o�E�4�ۇ�"��@�y�K�k��=7qQ�N3ʣ��dH���A����r1&�I��!�f��i�+v�cPh�H)"Ȃ��	�QD�þ��AWK���c��PeS��4S��_t=�M�i;�*w����YЕ�Y=�7�5ͮ���q�9��P�cK��籧�Sz�p�����[�0�Oh��2BKi*��<����ĥZ�@:>�1�B�?�`�O���_%�,��p^�<P8��K&���@��B*:̴��rȝ^ ��
�/I[��8�80$Ȣu�c�D�[+��#��7./`Ԡ�-�]��b������Ԁ���S޺v�����\p�5����[׳���.��O�?&"�o ��̡h������A�G!�
nZ��R�{�L�l\���`1�j�}���Y=�D�T��q��=^8�!�i�	�s�%�vw��$��<�P��bXlr��0(�t#4޾��v��3.�n#����-<�����[�����Pb�nL���j.���mgz�ĭK+�S����*���T����P��P/�������h�Hu�@�ۥ�%~�w��cB������f�iEm�g[��T0?pZ��o�-��߶��>l��*���pC荳�|�(6��O�[�13�"�+�e!r[�>�Q4z/�Tɍ�U�-�}�5E+��E��ա��r�+S���N� /�A(;� %Y���g�ٺ��K�Lp��4rG����. k�/�x<�S��/��vAw�=!?�Ql��!O8Ʈ��t���;���W�)3�4��3�ڵ#�C��q9I��®��`�Ec�Ӄ��X7Z����R�nɂ&i�g�f�"p1f��yMF�G�IN8B������T�����![�{N<��IC=2�B��(?E#]�>�o�V#)��Q<_A1�+S^@ND}�;���K>�m�#������Q���k1k'7%L���F"R{��"B�*���}-�}[�7�S�e���A{@�{uR(Ǭv�ޞ�[P#Y��|!$,����V̒�ˍؽ�(�醨�^��#o�]��3ّ#�{ԚGt�P��{����Cw�����h��q�2�U_���<c�i�UqyU8H!J�e���J3��e�_�������䊜�u��V73��U���0 r{����v���B��MM� ���/]��6"�p�-tT�g}/����jv��F���t�6ֿ���	{ﰘ"�&�ɩ��h�N~ZtO��g���kY�35��J�;�u�5��h�%�t�WU��Ɠ�W&R��D϶O����Ojx�֩M�td��U ��������xc��!���d��� 巍�������xS�m�S�����T:nN�$���i,ذ��
�u`YrpSG'��%��s͖�w��P��x�mZK��y+xL��İe�N���Y���%Y=o*� 8����)�1ƫ^zyӔ�M�������
O���]��	��_�+<��V�N�icw4������F����?p�l����[��_|�Q l��mO�n�#0���4!ç=Ef[O	;[��˭�<.&C���H�8%����xh��EZ?���h��g�Q+�����
ai8lu���p|ku-������ÛD�E�x�H��"��qNnm���?Zs�l��R�mF��	j)S����v'@��e"�5m��a]숢�>�ڄ���I']Xv����R�?�d䴈5�*�;��κ~D�� I�BWq-n���T8$���!��&3字Τ��#�w�R��.�K����Ϟ�U�/��}��3�D������<�������$��Y�sd?��)e��$N�؅��������)��=yV{"��4�������c�i��ߢ�T@B~�DjR鏧��@Ȱ���Y���G\%4S�<S��p����x}Q���,��߭����͞S�P)sl[%cvޭ�f=2�l��8x����|�nB�
��F��oZO�w��^�M�l����,��/v���wX1 g/:D8|�*4%/����	�y/�w`�w��\��W1�&�b��ʲ�XV*��{œQ�O���DX�g�d� �ּw��$��5�v�pS1���cI0��w�LL`��0�3��NexF�ҔA`x� ..�(8ޒ�����xt�����&�%3"����"=qݻ�<=�ӞvaZ���>��N{�װ�<�mq���^��B��5%:�,�9 ��J6��X�7u!�A��3O1�(ua����m0$5)?*�&�6���Vً\�"[a'���*�� �[Z#�q��{�ҿ��7 t�H�Ȉ�dr�w2D&��3 �λ��������jG݉�>�N�����X�3@��	(Y �������Yzk��D'�9.z�����D��`�Ua��I�"�{a.t::�@���C����R�+YyLӓ$�Ӆ�e����0{��X*e���t�����"����W����Zӻ������g#N�o�Y����J����۳���r�&����+����V�#�@�b�چe��Ŏ1��&oo3Y�����4�
�����,y��1|�͞F����s{��$�,�4
.uI�}G�?!���&�� G��n��Kޗ�[T��Ӻ@��*f�f+���CM��5���K���I:
�y���3�0�����`����^�r�P�+��ìU��foY���k+)�x��a@C�p��S��%�"�}~����#I��x)ًa1cR��k�@�zdg���s�rOR� �D4��h��('ڍ>��M.Y�E&m��rG�@d���@G�����i�{ٟ���PSXD�7�jD���(B<$,zB�{��yp�B��i�4��cFp#s�����Tʦ�Agq
�c�r�5��.���%�K�z%�ޖX����\�˪�[	��s`�������y�_��a��'7��.`����,y��qT�4�ni��X,$_9���N�=y�S?JNc�>��j��K���Pn�끿v�xD�W�wD���Э�پ��m�+C���<�*ݕ���q�n.��YX`�8�}2rH��D�:��T�2����OF�����?�N�V��k�v�* '��`[QQq�Dah�j���6�/��P��T�}�:Uۉ�|�X{!Q*���n� y;d���"�G�!��>j@�M$�0QM�h����5Օ{i�{���]���uS� kr.�����$�mc�#Tl��#@�T�� Q���e٢�R���V�<��d��G��{�Z��������Bb���gC(���n�� �/��t1"d�æ�E�A�<�E8�������a
$�rf�w��PQ/"��Q�<,Ϸ��siJ��(�r|�w]��>����|��a���/�NkX4Ə*֧���7��X"U.Cn@uQ֤"+w�Yx81X���Wu���uj��a�Cb?���L�����q�4ڬ-hx��~a����]lQĹΪԍ���w�Ug�8V�y$�@���;�%�Ծ&��nA�E�E���_g���~�O�3!�nbXCL1ov;��amH��7�� IH����(d=��\pu���)���I�����3����?1�yy&cF��֧fz(�Z�G��S4�1Gϭќ?�I��FW/,���Y�=Y�����%Q��%�NYT��gP�J{����z�Du&�<�t��j�� 3���L�Z`H��B�T�7���6j����Öd[�̽�91v�ܡ�*F�P�$O ��x�c�"��j|~��osO�5g$�0�/ʏE�j��;���sj�F]�ܞM�=V�����Z�
Ѩ��x�0����-o�V��0��$J"�YI���#��v@[T�&�Âz����`:N�FMX��fd?��;��܆d��`̗`cF�c�>6x��u�����6���n��,����	h��~�޹��M��aёݤ��;���;9YcH��N�q8���*�y��Al��R6DU���i�B�Qn�-1�B��U>!x���%����D8�c�[����(8�z�!U�#�����1������4gX|�����+~1���X�p�9
])VM�i���ɵZ���δK�O���m��f�'D6�lUn����mD�b �ܮ�HZ�jY�����ܧK�K����G�qg����fa	%�G�ª�j��K�����pJ^%��gq���m����_�1a�>���� ��)��Q���9������?n���he�GR��9����P}�H��(�c5���= �IL��b	~ _q��X��C%��
���G����
���r;���i:g��~�U���{���>��@�( |e���Z��BW;R��F���p�<~��ݙ'a]b�S'���;C!���xŚ�����I�]%�����0�U��Q!�|���������,&��G8��k���Ah�����^��4�z�	���f�Á�l���O�y߈�\�|����Ȳ�	��p����ݩ�i�
g1�;��e�2�8h�R͸E^�y�9��0�r&	�6�WvԢ	����9��e[�
�a���FW��㣭<k8i6���d{����"��D�}��k!�% �o`ߤy���2��׀S��S��7�|��>T���~1�;N�1s��D_�`�bm5V��LQg�9I�`�p�۝Do(����S?��{���k��c�Ş��}Hsc��ɀZ�NX���:��)�E��!�b��&�3�����8�:��m������Q�9s������&68�&i�b
��<if��i>p0��6��5��RcW�i!�s��U��vE��k��`q���J5�T��?9F� ��^Xq)T�6�Q��@�xB�y�hχ���w!	���ݘ�[�[���Ľ�%.r���nL�5wI_?f��-ݕ��+x��mi�����V�O=��E� EZ �L疤�G��|�~d����2��?[��m��C�M�n]�A�ʄc]��F�9r����=��;�h��~b�>��3���( ~�N�˓Y��G��d�<�� b�����a�n�5����r1K&ݮ)�e#G˜p!��V*�'�o�?�pg\�PЁ��.a�ޙ��Rg5j}M0��!�/Wg�F�k����&0*����n��P�*	�ɨN��:k�oX�-�"����?��.)�ʍ6� ]�I	��Z\��*�(4�h��f��inC!��=��I��K���������%�Ԟ�K���^����a�r���>�AZ�J����`C��sZ�Ǻ��6vI_�L���}��6�$P�����w��Ŧ*6E���!��$��^,8~EK_֖K���c�Ɇer�w-��L�u������a��Q��V�p�RD��8R�!W�8������E�J����V(��r�S��l!
����nvcBm��|���
 ��-Z�N�zu��%���$^�5
{Iр�����@A���`H�#�=�+��SGWW�m���׼^N!���0�]�;%����3|��:����������0ȶ���[��mi+�����C��e0�/���F�	�J;\��h5_�!��Ҿ�Hτ�95ĊFa~�-6hA��;��
�8��ws�d��'�l�ؚC4�x�<�!�����k3.��Āi_�$̸����6f����q�NpP�杽�Fؖ �,�@Al�%2L�C��5I.���Z�Qџ�;�H�G���ϯ��.h���s�Ƿۈ_Lp�J}B<8�	5��3[D̻��;��h���q�P�q���쮛�u�/����Ƒ��/��[����ׅ�X��$mw�K��@�wo�I�-�?�L	n����"��ϴ��l Ǟ��h�E��*�M�h3�;߆�q����bY���E1���F�=����XuYh��.v`�F2�Ŕd����<Ul����IO���Y���w.Nt@�ƬNP�K�u2��E�O^��`�~xݮ��2
u�Ԧ��<���ʐp	�ٳ>Y���!�Ӟ0�f�c�X<��З�\���u �PI���+��F���Ao��!)�ƛg�3ާ����D>��g�{��a],�%0�]QX1�EzZc�R�)�!� �ȥ��n)����������X�US<k~lӊ�;���;����$�����e��o`Z��@GH5*��&y\>�fRh�٣�{�5�����.�<�z4�/с՟j���7UhM��<5�k�����0K6��'���F	���O���_GF�!'-%e����2�q�����Q��.�6k�ʣtTA`VXVJ� 20n4D�r�^A�hi�z#ɣ�CC*m�$�*We�Q�i�p���}%��c��kT���ى� Xb�:{�}�ļD3{Nq߲�Rg��D�������tuNIv\��2�S�M�Aj �p�m������e��|`����Eb����Z�2d�/�Q���Z�w��N�"��W�8�=�N&8�4�:K�$�H�}k�����d�uK��8�U�KSk}���X�'H�`�Voݙ��J��x�U�O��_| ��W�z�#�q���
�a�!x�`��<�k݌��6�UD
���B	��H��#;R��[ae�~�ը�=fR�?�[���^��7�� O&F���r�!^ ��qP	T��p�5��J��E���a�ךK7v	:҂�@|d���z4>����s��MA�v�������,V_��k�??���\(���|�$��L���W~�S�n���Ue��c�i?��L����vn�bM�7"�b���0�k8-��Ǹ����T�^��g�Z\���V-��:
��M��9�w�E.��O��'$1�: 8�	B�#����:�A��#��	|T0Ǡk���'j��ܵ�3σ���Tԡ�
49�U��R&7�[���m0I��d��3#0�\�h�Xk晤������]z���Pc޹|����1l������>/{���{ި�-@�*���4�,l��Z���m, l�IϢT��+-���S��䂫���ߝtu �Jl��恗�T��6Z@��0~w�QO#!Aȧ�Z��nm(�O���ذ��f��K��Z:��Dm�[,c�dUR�.�����	��0��������V(D�h��!�BL�D����׮,oڏ������um�D/Ū�u�#�R�~}��/������P.w���d�^�g/%Ei�iD��Ȥ�35B�ʡC2L��,����/��<k?�I����j4����z�]�o2'o���DT�2M�()��{�/�sL�%�V�4j���<��zC8�.�#4���3�r��ۯ/f.r��&�k���0�,��C�gY|j� �~)#Ǟ-(�=Zy9Ly.�0��{6��K���{�A�Y&� �gB�k��ت�8o2����N&�����R�[���g��������z��c���r@�4t�<����((�G���nB�$�ݷ�*Nχɀ&)�x��F��/,F���X�c��,�%2/T�}�iB6ST���e����JB�>o��A�Q��̵�v�V����i3ͱ�C� �����2���W����3��6�8r98O���;�5�ǵ>f���L�����nwW�s�L�0�;�S�7�*������}�Ɣ����>��O�����K��m�}� a�>�R2ߓ�yM���v��-ˆ�Arg��(1�
����X���_&�?Z���j�t�ĳⳌ��Z�b�5�FY4A��uр)^=F��kŶ�k���v�݃���[#����˦�j��fe3v�*������%�Q,4�K(�j���q��S�)�jUb+�b�g��w����v�l}�6J�˟���O�?��'��h���.~��a�Vr�^g�yM�?Ж71�a3Z��7�]*8K�*�qmt�B����d�6���*qV��8jpIྸ/Q�RP�!�#�:�2�}�r��p&QcM\�xޟ2�;���W�p�Ef�c��[��!�%'�%���P�<YE�A�Uz���V��"EHa�(x���7D��_����6[��{3��-�m l���ar��5�6^�&e�2�L�E";!��0w�8,�44j��`7"$���1��?�w�#��~6F�X0!�~�)����M�P�쫵-#-���Oe�GLzb1V��G�#E&>K�AR~͹fء�@�.�$��)f�̬b��x��%����b��q�).fMulSC�{J�xW���0�VK]F6�ހ�s�l����s���/�e[f�6F�|����P��?��G}}3v���L�3�Wk�A+�����q����w�_�m�͊�Z�*�i�KN�Q�])<n�畯>��
v�_�lw�"�c�w� �������o�<y��l������!�����v��4��^/�r�H/�a� ��\����`�DQ�@��݄ѮWJb)��f���7�r�p���g>H��!�_6�-�4)T{��
S�h��e�t��'���/�σ��YA2p�$��DU���|0�6�@9��������ns�~�L����<���3�\"x*��šS�d���]��'(���$/>0xЪT'b?�". x�2{g��!��a;�lK�`~.\$Dk�ǟ����Pc���?m���e�md�����|�ʁ�U��vUJ��4O����a��,7��n�S�a���`rM=!�qn�D�o[E�x��d�0Lk��%)ׇZ�	��(��R�%�Ӛ۾4B�[B��U47	�&[�T��YG����m�ƭ���47W�x�;>j���$K��;K�y�&nM]l�C�Ύw�Q������J�Z���<�����E�1z'�AN�Ѽ��\���h��6/|�s��ęVx���G�$WʰD�%M�5�����ڱG��f,���+q6M�R�.�����2���<��%�} ��?ܓu�����P��\���wj���'��Bė��9�Se�U\2����/s���Թ�{�0�\r�rx����!A��@�Q����01�+ފ(�N	����dn���?ٷ`e�89@�N��i��f�\v����mmM3Ā�+>�ݳ^c�F�.P8¥�]ϼk;K�T3s=G�J6�Q!���q5{u$��D�v�r2�P""{��+���C�4+�ˮ���29������`<,3�[�ʁ
a���H�	yA�2S{<g?}0��4��z�� �T+�Fb�-g�J��3X-��7&��<\&���|��\m���\�ܷ%�Y>}����1	1�����_-"�]m�����D�o��M`���z���4?�("*(� GI��/}��1y����`�f�Rx��V2,A����9*�~�\�J^�jy������5MًV�[/%q	�:��<�%Do9���Yq���ΰXC A2b(�@��2��3�aV��?��m����@Ē�L�Kә'~/�U�7|4��.j���5����>k+4H��U��u�&��9u�檀�����5���f��L�,�牄�C�>����&��F3�u���w�n�F��K�3DL��F�_^�b���1>S�9���<�oF'R�����9�u�̫��������x$��&6 �SM	��t�_
�_�1�-j`\v2�u��m�<o9�ݍ��к��z���Jmk����h�qξу�����-P�q�;�(��rQ���6�w�VmK��qr]gD6oҮ9Q��;C���%C ���
w�����s�
'���<���v�{�x5jN(Ճ)V���
̺-Lu��y��6η����X�fa���.7�i��ܕ���r��tN���X�N7.ͻ	����zyF~�z�i9F����ʴ�|��˿�d0R+��C�#Wۘ ܧ|�ԥxp�v���`�~p�Q�
���"�Շ�|��ǎjBg�6H`
s�Qx��P)�Ti,bb�c�P�%�PX�]�
#�w�ԉ��d&������6-<�k�{jo��?ew�D�����F�h�P=~�O6ޜ����u}�6gWl�Q�?>W%=�������f5TSvٜ��LM��`S��ڛuX�hw�\�Lymq�f���/�}ʥ��v7Qmӫ�W���һ(-O��Hj��n8�9��@�%k*"���"֑m�1�^}ٍ�`��00�r���U�1�
���}^u�V�k���畎�x9�s��-�%=#�d�	������s�@R3z�aK�'�\�L��0�O$�;}w���~�!Q�\�S�`Z0N!=1��(���˖+ډ`���0�/�����-K���$-y"r.���!+���+ R}l���ʠ�
{���ū�ZP’(͙+��2�0�-V��(
��! p�rs|5��ӆk^�yMRkĻ�o�8KR{J�7���Φ@M�F��BU�si0B+�rW�V���:ٸ7��Lk+L�̆5N���h�]����Ρ�|��	���2>�W&��%��r$�_�o�7��&����o���v����X�F�����X���@Ȼ3f.r<E�*�6���׆����TD��Ѳ抦J��l�{RR{<
9���� s��42�bs���o,�=O�f!����rn��_D� ����, ,ϋ�5��1�#���@-f?JS8;a;�<���Ύu%��F�[;m���L�%S�9 u�u���~-<��5Y1=`�(C����8��s@��� Y"�m`ɎYMQq�p��Î�L�	��A����O�4r��%�6Y�u���P��g�2�.����4i�����,R��S5m������Yz�ݲRo�eD azά�%Bd��s㞗�c\`��K�Y�����!�hFkn<<��(Hv�A���a�V`"j�k��5E3�鈲��᠃e y�՜f���n�܍�_uvn�y~�\Y���[�ȟ!)n���bN��"{�8u�+CS��ᩗx/� �RJ���r�F�J�rK�B��jrjA�	��}��<� ���l�^�S�IM����Q%kV�"���-G��ƾ_޶�����:us�Q���w�.F�~cQ�ɷ�s����^\�ϩ��\9��r��EXmDV��B��	��5��q9��@���o���.Uz.�;1�'�dnw�"G@:��
=uwb�.��5��~1�w��a2* ^:�CLI���L���Q	�w�ƶzQ�hR�'6��!~��Ù�-��ѿ\��a�Cd�fc��0��DHqP�x�&B-%�ht�n\!w�k��8���)\_�#0'���˯K��g���Xۼ%��Ȏ>+Jt�,���Hl̹�4�)�W�b�ŮJu�R�U��u[b�o��d)Q��Ҟ $�p�yMY7���b$'�'��n����Ʋ$D�8�H��o/I"t`r�8v�&�x�⬂��K)cj! l�;���Y����w�����XmXy#� ep��!z��MF`Ͳ'@
���f��ʟO=&A�(� �Q�S�Ӫk�Ekq�e��H�u�j�>����k��'=�ٴx��&V0��Twdt���^Ǜ7+$���,��gm �=�?��h��Y�5��mV_�?B���̗�v� )��W{y�b��me*���F ��>F���z�6j��3�O�YpF���8�݄앁�m�/1�C/���9k�MdI�o�6|x	\S�>@�x�񁃕O��q؞Z^ؿ�������Me�B�Y�!F�9Qa�ۃt�q"X'Q���"	��X 5\V
��f�B{ITBW� �j�x�B���_��X3�����f�6�u�����%�.������{����b�z�c��H�*|HOYs*�g�P���dG�@��V�����l�=���-��U� ���ԩ�[X���Msjh�ǖG�P�T���J�m�R6]U���C9�v�'��ε�9�2�ȼ��a��Mh:�VЯ�)*8�r$��o�e�Sr�&�>���Y��v+>и.����RU����j�d�ϻ���܍�?���z%�#��u�S-�C6�b��Y����TB�P�I~�h�T�j����A}�B?.������^L~U[f0x)�@+��?�h�Z1}�L�|`�ޓ[= ��Y�uC�*i����i���k�b�L�#�� j/��0(�:����ۈ�WųS5h;�-:��eQ{ӇNU��%<J��Z=�Vd(�����r`��O��z(���PMl��I��l���Pte�\R0�>�IC�>ӫ����@
�q�7rD"�ߖw�Q�S�˂����	��Dc돤;�g]i���|-Qw!�(x� ���h��o�_"8&� �vR�
��u���~`���ֶ余�H��cb��h��$���7�,+*�\`-��ܶȩ���fA�'Q�y���d�?�K����щ��Z�+7��I���[M�#-�ו[��Ke�otOS��.�[��'��lfVnp���G̯�>��D̷�o��a�E|���It�>�m�}��~�U$������cC��MB (��Å�W���,��б%�@��������%�3�9xP"�SLx2���}5�`��"0�?�X-ؑIn�n�KԾ��D����~�.��rV�*�QC��;W	=� n6P ��R 	l9IR阈k��*#4�rǼ�Y=��:����1,�zsxiZ)gXFԅ{6�u&�#Zi�[qW>�,1~����������h^��ԋ�7ě:W>��=P Y���S<��z>�p���MU�G�
����&�Ԕ�N9���vx@h�%9���̦��HǮ�'�B`�֫��{��b�hwf�j��On�����������H���<����oi���d V��8���(n�����Y�B�0���y�
�/��+66�
;Du�% )w�ɍ��J]N�oj��m�b�:�[���5���ع���h��}*�8�k��"`���Q����J|]��N�^�D��p}��� ��!�ޡf_� ;��'6��O ɌQі��x�ڥ<��1���P���`�c�l�2f�'c�%O>���t�̌���J�G��Xsi����f����cU�5Ъ���_�Bk)8���n�1ER���)!�a K7=�[��T�v|�����Q������`O��8 �xg�$f04�F�v���ic��W)%�·�>�{���,d_�I�,��PH���;�)�">�3T0	cp��Z��-E��(�K�kje<s��U�Nb`��&]!.v��9v��V��x\��ԣf��]sz=�-ݥ6�f;���^�h����.\3����eu�j$��(��Hk��PD8%='�l/H,��H\�k[�e�S�g���W�/?�i%���>eu���y[�BL���_xc��6f����v>�ES�U��9DG�s�֛Kv�:�����'��«���"S�3.�b����n��m�������vjY�'}{� lg�o<GE�����r}�-NCʪ�\e�0~P	�]P�2���^pwz��x`��6��E5�_jǗ7I�M�o]��e�*�̋im�4~(�B���	����ђC��L�҉�e���0<��cՌ� H8Y��?׫xZ�#L:�W�g�&̭�_}�&�A����}]v*c��%vc����^$X�M7�T:Qf�آ�/}:m$��{���}D�Y��/S��ǟ����p?�a
�6Z�����W�|�W�sۀgT�Ӂ�8o��Vb��u�����-Y���@g�z��:�\�.�킵�	��@�J�؎�h��?�&��y�p/PҏŞĜ�s���#��Xl��y��F5���um��������T�����y|�{�W�z�K7�	�9K��8���o��C��
Ç��|�
�]�r*�Zz}FÆEoN,5jc<�	}�����h��b`\���S�z�N�R5jV�l��R�N���rh�6*�����
�7o�R�������^��?�"�w��d���nX�I��?�}�E�R�-J- � ��3�cɊ�������&Ӻ{�1c�%�Qs��>�S�G�v��}�~GBj.�J�(���ܯrzC/$�[�����֋{D������$2/�<m�U|j~a������_+Z���p�6K^`��B�"���U�v�����A�"�_�sN�+kO�Z5�����MOb�����t�v���z�����J�����<˅&�!���^G���V�����?Q�Ǝ-,���~9nTfʡ^ ?K����<@xrd)藢n΃a��ԥ�����b�Z�O\Vtˠ^z��eq|�ڍ碒�v��S��|�� �8��	��y�5A`ěН����Lx��,�F�b���jN�.����a孝�K�*P�P�I��� �7KDu�j�l��y��ia��(�
њO�:Ű�}����@.��!�?�C�@����Z�_�ŕкia��]��X�;��۬�czG���1N��c��@�w��տO�+��bӓ��Y���'%��θ�6��Ɠ���Bl�Tϰ?�ed?�GtjJ��$�^�x)K�I~J����F!��oJ�9���Z�T�r}�	�Bkԥ�/�{��p#^�@����k�NM�oM{v��ã,�W��cɲ��`h�#=�.�q,����O�Ŗ��kZB�,��_��u����V`N$w�'w�D���~^j�y�>wyׇաG6�}��TC �A�l7"�3�ؾs��R��&!��L�B3Xu�݉f�E�k���*$�fz��2k��)I�Za�g��8h��a�������<2x���t������1�ˀ�
E����|ؓ��"Y_��<��e����(�&���߹d;���=<������h�˓��� �2�{�"I���.�)`�|N��×F�j��G�.�����d�������O�d#��>xL;�'ҭ�c ew<���"��H��O����U�����{$�,�s�1*��o�Ğ��D@�Xvi���|c"TdrRӑ����?<^$�R�@��4(���B�,Uy��J�@M]#R�?��c:x�Y`y�@�71��(OB�ӈT���u�/3E]엀(?L�5/+��cU�F ���y�|������u4`P�����L0��PrĜ�1]K	
y�S�*e�<s��9�]��A�[�%Y|�jg <hC�=��OӚ2��	�C&�ʹ�'n�X���a�o�C��6 �5�)�48�yٽ{b����[��?6V6~E{)�r��yl(��JSo���eːg�'�S��&��[�G@��]���:P��"��z������ˈ�r��T���x!p��i��qy�9��-�&��R&�M`����T�[���p���M���O���X/�_QhM�<�#B\"}�:ZU#y^ �Ǖ�K�E�Jv��ċW�%�66������P~I0Pg�O~P���qiTK�0�h0|����BGHy�f�U<.����y�24�.��C$�	b�[�͝�	�th2�iJ��@��1�MB濭3edn�`��,�f��)�C�߬��S)k�%TG�z��0���'�9�/`�����=�9���9,�8�a�-�J�@�J��N�V iq_�]� �0(�.�N3�}j:���G�pȵ��.����.=A^��~M�<P�a(��V��\#m���-�a�P��|\]Ò�o�*^ʝJ�(V�9�U�����@�d��Wkl��|��H����R	��#dh��U���Su[P��'���'(�C�[]a�>/��A,����J��K�y��I߱LY��j������:nO�&x��F4>Xڭ$�+��7W���8W'���<h;�k�lJ�b�"ٽ�NW�ݮ�)��W`���;�QT�u�iM.K@�s�'�y��6�l'������Ѹ*�OEIC���:��
�v�]jNܑ�Y�S��W�
wE5K���3�1��k��;��c����gj!�<�}�g���sY�\����D��!J􃘧��t@��z�膾�VO���q�.�] ��7��a�m���˘���C�������-����� n�h9�\�&���<	����~)F�tO�b�E�P�F�AU�|�X�I�ێ�b`Ä�K̲N�9���.G'Q� AP8��`�}ޤې��5+��`��܌���{�I��5)8����@}�R���_�^JA���g�X<��oE�h��s��{S	zn�R�^+f�W�?��`q��Ǿ��`DP�$%���ф.�װ�CK%����b^z�g�(��GW����l���KS/vڨ����Z�qpH�UG3�!<�����O>��l�[㶁6c�h=k;�z��gta�V��T�Kz�	�#z��W)��MY����7XטF�S)[����铞�c8���{�5Y�7��Ty�x���٬�Q��1��|iQf�K�B���4�ń�rk_���:�^<��Xx�� ���d�J	{�p/��ku�.�ӷ�J���MǪFhv4ߩ�J�(�tv�p.6��D�e@,���֍��z��e9�OBX�OVQ��Xi�7�;�)����Uj�NJѼb���Q@��,0��|��O@��)����=nm9��z���>�#�2̈�j�¡n�tN��#�mef]�dh�쉴�/�H+/����&�vw�|��r �I��N�d��$&�]��+�4{-�qm3���N��Z� ٢R,/�vZ�.l=�t:}�w:i=�8x�;�F�Zp��  �XL���*�2��ϼ�]������\W	!Ѻm�cxY�]��G�d"o��L	T��l���r���Fn|�-@�W��[u�4v�4��z�_HTy���0󬊾��I�N��-˧t-�Q׮}�h�!�m��c����ya�2M���[�����wm�v�58؍�h�SG��3�R�-}��*Hcܗ�En��`��:�k�.l�l�����񗨨�$V���<I��ބ�7��t���`4�J�~Z�+ZOP.e�Zo���~潡��g���NTP	��ŵL���x��qUn�8:*�������@J� C�Ã����V�I����NMB�mF��O��U�x-�.SO֊61��{a+m��`g�8�����4�>nr��I�5�G笍�#�Rꛎ�4�w��:�ڦ�z�g���I��E
~���%6��%�!vG.�4��3;����V(9E,�vҪ	� �C����f5���w%����vhm�O�6��	���e�I��+K6�ʟ4!'lF�9��S�v1y`����r�mzx'���Ϗ0u�[��֣�bS�+����*�>�}3M�r�Sþ��d��h�,R�zu���=�RG�zV�:��'bo=���Cރ�y��Mtܯ��}��b�[��s�q���|�1���a���(ċX�����B������,�"]0�ٱ�M�S���$�i]9V���G���RF������	M��͋����Ŵ�P�
;��Ւ��N1O�%�t�:���n���\�����-��J�:�A
�� ��H�Z�v�ѩ�p�� �5dU�5�t����s8eht.�c*�i��J��c	 ��x=��:����`�N1�����=A_;<��6���B�������]%#������)���i0J�j����hP�U.�iW��+͏���`�ÿ�+��`���=pY�{�&�p{����+GCy^�j+��Xae�	1�.��%_�BP�ˍ8����o ���qFQq&�2Ц����w<#�Ѷ�,�2��EN`�/I�����ܼ�N�+3��K��v�qU�)�w֠���y���#67K7��1��L��d�S�����hl~4´`�-ҹ�Ӌ���bPp���D�H(A��QK�_��-GZ�"�� ��啃�D��ZH�?EY����ٯ�<`M�vX��-{O�hIϨjd�Y�iT�(9�IʑY�tA�p/���nW�t+�v��g�^
���x؛m9��` �;���b�&�:¥�ki�iy/�0&Wj�d�@|xoY+�"��L��t�E���	�jB�Sm��^o�>!Ez���kF���q���Ө��Gd�-��"`g���J����yO�/���ǫ8J�;�g�F"�K��G��neI�����V��k1C�"�}�YժA�3�^�9��1���3?���FN�Wj�#P��lgz `���{�@X��#0~'�0y�I�A�K6��ς��؏��pDZui|cD%O*s~b E*8zG~n�+�0(v!�Tk�+����4��k8(=o<#�;7�"�\YeJ�1u����ϻ�� ��[���\����ˍ���D����K���Q����d��bX���+~Ľ���ZBۨ�/<<UoH���MsT�S��Kz� !����C�ټe��ƭ$���
>��z���I�DXu	��O��i])m i�����p�\�6��M��m0S-Q9����]�B�aX���T�`���6��mm<y�����'ad��"묲J����)�W��+<�����H|3�dF�:��wZ����vܨ�CKUgF��E'(U)*��0l���oT�&7��l�Hw�����5��Rb�`xlG
n�"���~����	q�d���v�}���N�	�ȩ>�}��]�H���\g�x�RU#�%���W�)a�ȁ�7��:C�s�����9���@�}�G�f��@��.�{*������Vc �{��4LJ��$TA��)ݞK����jI��P���H8�����2�u�����.Щ�(��7�M���@�<�:X�cv[U��Ǻ,�6�2F2�9�|$&��x�`K�0���P�M!{�A8?_e�� X����4����lϣ��������*�e�-(x���K�)����ldl��Hà��o_�9�X~л�l��;M�:�O:e2��Dz���VP���:��>�����SA/�A�%�zq��c��;c�$�qR�A�Pۋ����%;x�� ��|�`�@��JO�i�4b�e;�B�� �b�|�t2^}���Ui�d�'�F�#q����p���Y�x���oj�
�+U.\���=�	{����I�Pxb|9��$gX�3�;���DUI�N�RC^%��
��^��.V]g�ЇC����_P�ԚQ��u>�پ8ng�w�Q����]-��}d��8�D�'�`������!�΀b�q��g�����?������BOofS���b���U"��o���M*���ԙ�����K�h~\�IWMX��@��GB�K�e���.�כh�Bɨ��+Ň�:_ª�۲Ωl��c����,�2r{/�ks6���`w��BS��泪�A	7t�'L䝬0�ůJ�!�']({ye�ztc�#��`�~�`{�Aҏ�E艘�A�pB�RsO�ҬD����B�4�7��ݥ�6w�~��ptȺ�ߨ?]�彰@�	�;[@������V���J�c6�q��p)�w!W=hέ�5�;n�Zz`,˽�Gpz�.�uR��;6�����?ro������Փg�31��M7�<RqP��	���lQ�g�T� f��O[���=A �?�t �O�x��A����L�#���`�K��ั���O��+{�(�1;�8�e�]C�ҵ�N�'R�C	���)�.C�;��h<�&�3��!����!	K�8���Go=I�u7�Ѧs�1����\�����+�Q\��M���l�,��sJ�Z�x�i��X^=���ph����w�)o�+���Q�H\�=��Ijt]�S���%CӃ����Z����b�"pC6y=��o.�O
�=5s"�G��mD�į��/7�����d#�
iʗS|gSS~
����A0W�0l�.||[O}�j��c�.�
d�7wq���6!e�+��زqb�w�u��y�ft������=b�`&��h~P��f�s-O���Y��b~��:W<�;
��܃n�>_��k����R*U��U"�}��٩F�nƈ�C,�L�[�vz&o1u�A�����b�`��.�EW�)��\�ǦȾ�Yp��*<��$@0}d&�(	�¯��Sg��4�|Ŝ���zg�ޯ����J��V?��n�Р�ap��T5E����ۄ�{~�|"���:��5
�0$�=�4�o��=��R�|�XW[�+iA-�7���A��UOB�5=rkŔ��D�d8j=�W��\��2�BZ:���LR4BdL�x�1)E=V��k0Sט���2<�V�u��G_eꘕQTE�\78WB�502	�dkB���\E��-�b��Dy����|]��읐}Lw_�	EOG~��h#��h�V�g��qU���ՙ�*=�{/��� ǐ�i&��K�%1�z;]j?p�.e�wBx\~$M�Ք58nds��.�a��ͻ��Fۡ�J�Y�V�� Y��JR�f8+�͕ }z^!`IbqOy��(~3S##�h-'�#`U�L�	�������f'i�vLN,?��z�M�2&�L�����iMq����3m���}�+�"z�s_C:���q�d��8�$�mԣ(-�k���ƒ�:0��I7�FH��n�j��S�&�콥 �m�ȱr��yLL�X�ۂD1р�[(�I����+�%b������abjRX�3aD���)Z?H�!|�ۦI؇\p��Q�?��� �P�J�	sٚ2c/m���:��xk�^Q�p1i2$��$zs��t� ��Ee1�([�ӿ?�Mpl}9��>?�b<
^�o��9MnƩEH9��".#�5uŲ:B)����9\��ܼ�#ީj1�n'�n�m&z~�[`1�܇�ge V��[�E�w�fD
!ޗ�#R���
�_�vE����j�n�0��3I�P�lDc�ӿ?�ܾ�i�Ic�:����DDo̔����,�Hs:��j_c�c���nb��k���4 㧇"��76ȵS��e�Z�rr�3B�G�m������`�_X���a��|�`������R��z�/;U%6�^�"�Uw.�F�] ���b�=�<}1s�T���dZ�;��rl��@	e����Լft{��FL#�b�g�V�V���	�ie�2���m-��L�^����VJ�A(2��X���f���&L<����_�M曊4%�,���;WAT���%�OL�t�u�=��z��Ux��Yʯ�l��{v*�{����������S��fln`�F����9��fCh6��\��N9<�\��!xc���T�z�R��V��ɤ�_�3gǕ%�CI�x=����YN�,���0R��%lt�Τ�@V���9*f���3e��������ڒGkO����#�ٰ$�ێB�����&�|}���~�U/��-OS�&����cފawM�x�,v�a톅����D��Ց�U�a�'@�d���R$U�RJ����TV���
�=
�>T�2�� :gh�oE4|�o�&����>��u5)�o�GO��M6��g{����������|�����l��Ep��!��ԣĦR���TW�_�Ͽ�"��Jݤ��P�%.��g��&�pq�/�Z�6cS�ލ��.�񯡙�.lݰD�K�����%��1}�b�܄�D4L�:����ꌱ�� �pr�T�V*�1��Y��+ϥ��i(\>��ne�D&:�����spMD�����I+UU�ĐcGX��P�Q;�~aU��k�s���uf�H�w�vmc�O�}���4F�m�^�OA��)=[��4���>՘q3(�u�{�{��g�Өl����f�J����I`�P �j]�.r�1�]���MHy6++b3�'T��[��)��~ST˧V�m��U��6��"#I���)m@;�nՇ�%��彐�G�ùmqRT�"�FM��a���t�� \��{��M��ϙ����b���=Ŵ��
)�������	7��Aw��s8�U쐆Y��|"�����ĶQ����Y��I3sl\�B��or�J��-W��X�MW��7��(�:L�5��p��4�t�kej= ��8��n�Z�lg���$wWX_�p�S=,YG^lН��Qş ��V
~d
'��z�%�y$�6���q��.���_+6�ŒZ
9���l$?�H�a��KRޠ\ō����-�/��,�ś�Y�n�O�ۆxi�hp���|�ED��g^ �"���(�Ϲb`�+���d �Ȩ%Q��l:�W��C��]͌�<���9>��>�)DQ ᣙҗ(��F*ۆ}s�<��A&����H
�� ��
�@2�S���8�R�
�ۉ���>)x�ߛ\"�����I�Y�,��ז ��\��?}ޗ-;XP+�E�*�D aԦ~NX��舗 T�Q5�h	�\��P���Mr���⹱�ɠ	�W9j����R�W��撠r���O�w����l��rg=0���'WWDJS@K\���B>�1�)�����%N�ln���-�e�y\�e��e������9d�������~
e���gǍ��hH�Ķ����3�J$쳐���_��f��r^	��	B�l\�.��&�ޒhV�X�<���~��z�/%����k\7ӈ�mr{rH�➥,�-,'k���h��~�I�כخ����*eޘZ/���Ľ͏ͫp�ȑ2�u1�oy$��)�]��)y+��?eC����i��P��1)��4�	5Iʾ@�ּ�5�!0�E&�,�U�i�k��%\�rDs�OІ�&>8ݍr���Y���󢴩��=X��0�YI,^I��l�?4�ב��3���-�~~����r����Ėo�|x8C��?6 ��W$�y�\�̮#���!����!�����3qE�5��p� l�R�Sa���!����ǌ��;�Z��͏�������?U�|���������x�#�G�y͙ ���d��nY��aQ|��8޵��ܜ�gj�^w�him�>$��̡V�<�:�_�W5F�2������=�L+�x-�c5-����,xl�O��4xfH���ݼ�w;�5F\�'+�'#���yP��Q�u��>���c5�U�ԁ�jN�uL��:ٰ���+�!�\�G��~|d3��#1ʍͫӊ9T���2S!q�ߺ�٤�ֻx��ߒ��>W��z)[��u��h�WL�~��Ɂאuvm���zh<r�Co7��0�,M��Oޢ�{�Y
�yN,-���y�ƛxF.Aec(�Ah]�#���a�8Z�I���1YUZT�DG�4��`B�"��琦=^����eG}���m+��1�xA�Q�U���S�W�?��H�u3�b?_\a^�{(�G�n���|c�K��������-�T�R���K�]WaumCs�oC�;+MQh�9ș���A� ���W�=�_�����+K�`譱G{X7�-���\�q�NW���/`U�[��������Qiw���'�\�^����A��Ѩ��n �94]��cI�&��<qqD���X��|[�GE`	���A�oj��Z	���ŀ�#�E=!�YX57��Wo��
yg�&:�2	��-��_��Ǹ'q��`S�1ke�n&~��M�ceB�������>�� U�����`H��&��|����%C��3�f�b1���q��"<#FC�*�ja�mY�H=F ��_�R��p<�8|P��t�B\4bì@�@H���x_V� Tm�S�++e �2�'����F�$,Q���&�J��F��g�?uS��(�L�D�^�>�"s�x�]Fb�����	��
��3�]�`s�)�Y����xss>ݵ�6���
"�#3����[cYⵙU�R�ԇ��MzV�T3�d��P�ݤ�m�G�xݼ���Kµ�7J5�YP�3�ɀ�E[��3�2�ϳ������=�R,���6#����c�&[�����X��<gB	'��O�l����.�d'��K�~�A��,)l��b;�
���%'+׀��Ҭ�t���$^��I��k���sZ/��'�$lcqn	eK�ƈ��	<)���|�W,lj\�}�]ߩذ�5/#$��w�L�+�K�Dz�D�L����罹�;�Q]P���+7�B��=P��8X�gL���8MJ�K�=;�t(�:�l�������/�a�����荥Hr\���m�1��~L�l��i�'ՙ\]m���۾���P���[����گ�v�)6����f��j_;Ѫ��-=)�^R��!;�=�#��B�Ҭ�)���l�E0 ��7�ԛ�`���_�O+)m�]#O�k>�7VE#��'*�x� ����1S��(�B�B.�܋-���A�CӀX��(h a��p������mj�>��b�m�a�)��
|�p/=p]VB<	�7�ލM�8-BYob�Y�#EԄ�P���3��x\b6�V�M���z5jI��Q�����v��"�Z��|�㣖A�>�#����*Y5|S\x�7�bw���L�X�)��/5��2�=�"d՝F\�}��ˉ:����>�o���G3cb�b���2�UP�]����T�E[�M�ywF�81l��m�R��	5�#y�e����C�*��>'���K#͔������L;��cE�+c�F��3E�UX������(+z���	3�� c�5�><�M�u1,P����"���H�<��wA-� �v���'�V5D�g2��j�A��,[��Ƌ�q�q@,�eН��e�kt��	"R$nP�HU�e�}cϙ�������o5�����Z�R����R�6,���[�ǫ�J[y,�{�5���W!�~�f����y���!�I��/EE��a�0�� |5�<fQ#�;�)s歷�R [U_TX�`���U��%IN�I!G>/��3P�{)���<�|��Ղܵ�I[�	:P�)��J{3U�T��7!��̫ȼ4�	TA�r��U�ȮCg@�@�N�0A8��/�-tQ��Yf?@�	c	2��;�V�\h�g-�j�FG#�Ł%~�P�����j���m�|?��=\��9�H$f/�)Ey�%�G�.�J�xs��6��{v�>,�;���8��f%��$�Q7H��f �)W����J�K��߳(�Ǆ�Be����V:Eo]�p���֫7?:��-�1�(�V|/YE��\�<�l��+鈱�y)}�>A�4�. WH'7��p6�ܱ)9t���������ߘ��0O�a`|9z��A@=7�L���{4B�R�"������A�'��^M�)AޔR$���w��O��
��B'�R���T�W}%z���!��=�K��FAɋ��\I�s�`9�v�5�E#0St� x�%FϪt�Џ�����%��"k-�=N\ n���t]��S�.Bi�BB��G��jR?���N�iE���0�	$"�{��6ڒ���d�|O���t)e�zC��$�>��0(L��8��lo�rc�3��l��G֟����&(R�(y#������3�o0v��a(09�*���Qy%rԊ}��@"d���n�+���:.b���9ӚaQH�2 K�e���D�k=x�yn���
,��j�$T�ߩ����2�"1�(�0# ��!�;��^�sܩ�#!v��X���^�^j���{Y�� (�x���W5y�8��"�3{:�(D��h��6�b��� H�X�}EIo"\6�֍��vV�S�INg7C���)���X��l�۽��p$�{��#K������e|tb9�W�T"YJ����_�W��3ߙ$dp�܏1DN��\��pFQǓ�ɀ(��Ě�$Y�V#Z�YX\"N_�����p�Cq�����kS�ĺu$��	�m�n�;3��H_�Q���\�H�ط�!pm6ж��K�Ҩ��T�Y�34���wU�K(��MiӶyI)"4
�m�˳2J�ml�9|��-�e��-�9�fa�=��}���Bh�q�	'��2�@��;{v�1ۺ{�~?B����c5Gۨ+�>�{��h�930%��H���O�t(��h��l�x�U�Hq��5S��3\*���m4�<�
��x���	����p�t�!l�\�:fB-G�¶��X�B�䤕p�fK���<�tN���-(����ſOBT�7#I}�N�)��֠C�V\.��U�\t�YިdϜ��V�GH�cI���js��@o��h���!�r��}.��*s�V�������)�绬z��R|�릜���ҁ�=3^a>)�G|b,�
-�Ft�ej���$���lьC�K�$5>�����	�q�0�t��j��s�(	(�|B��Էh:��>��*J�L���(�c��% ��([���XV�Y�q�/����d���s���.��qaBWZab�m~:O����A0E��O�'b�C����f���)T4�[vn؎�o��$��E7iDx���&�WU��%�r��M�#���;.9���	^��TJ���7*�,���T���(�ˀ�	���ʞ�L�����u{wh�ώFD����UWԒW3���I�b�t����&'��ޗ"J��  ��E1���F��vP�E�Z=*�_{I�
��ZJ�uz�'zk���r7�~S�y��^�R�T���(�WI4�`˾���/�������5.�m1u����i�߰׫�Υ�.�irl��\rp��5ݽ�'k��0]�j��>�k6���u0�����=[�l���c��_�i!>h/:uI�Z� ��R���e<"�&r-�Q2Z+�U6ϿC��;(�2sd�̔�����QE+S��`K����/&K��6`��0$I����E
ujB�t�{;`�o<!'�:�=�ܣ�p:�n��5�Avlv/��w�b�o~���B��Y�w���mފ4?��!ON��w�d�)B��;V����}��+�1E��\�-��V��ۦS@��F�X�����ƃǞ��}�ds��n,��ϴG�g�_H9����ه���w]b�UH9����?@�� ��(Vr��kz��{��ު��W{Sa��*��_Yz���9kM�\��\�s"F��b���!t�'`sw�ҳwjU�w��'��t#ۉWL�B7��ègD�3�e�>p�ty�dtw���wI����e�����u��X��V{���nO���C��߳�&��K���/L�:��h+������ʐc��a��Ô�Ϯ�02��j�.���6�� 2�_���=n, ��lU"f=ʐ�n�z�|T����GƞkL�z?{��,i�ui�Xf]�S!)��3K51�q�D�s��i�SL��&;V�$޷i��h�`C�:Y�����ALJr�� ��m`-~�P0&��ԜCϾ`�:{���H:�7��I�x�%GC�D���������#�WĜF۸�ř�&�{��)�t��Jb*!� �}�B4"��E����s���<��S�y�w���G��^���(��>����o�iz�b!��\�t���Y}X��w��Gt�P^ZuN��( �:j0��h�Էְi�I��Cob�~�^��x�!~NX��[c�_Ⱦ�oT�Dl<�1+˺��M,�-LX�֔�F��*�ݤ�.��4T��\5X���{^8�V�t�3X.`7ja(uW��.��)f����.����r��;��tP4�(*{[?��ۭ�����!���f�Xh)��;I�/����h�$�۝�U&�BfB=j��:"^"-�`���|%�~���uX9@9���Νc���܇�/I`s���p�ݻ
�7A�D2B��O�7Z�;�bXi��@R
���ѵ�U��폛FW���)Gj��H�IyT ��
����h���H͑��vY�~�?�<g�{������_��L�G�c�$d�T�)-M-��V�@J4_0y��W���99�Q=�{�p!���F�!oIm<�0`�����ǽV�D�#Rd��OQގ�o�L�R�,	�1p�lz�ׅ(E�?��?D�[lg�,d��5
�䅨X����G2� ��=tid��|)���ͩ�ţ�U5��
��]h��0� ��&,I)Mƪ�䇿s����bVI9$����$x��k�v��*��܂�_��c�c��D��y�*��(7���˷������o�������%O2�6�������Jw^������f�z-�"��ϾD�;ܷ��_q�gq��c���$K��ԛ��'��~�#�P=$z	Q2��Տ{eRso�qRd$cw6>���+���4�E@p~���n*�C	�s� ̱�w��I�Q�*��w��{z!�θ�P��=�`�C:�O%�c��KmG���N����=z�ʼܹX)ۗ#�f�z0��?Ȗ���-aۀY���lyy�ҕ�"l�⧂��H2&�C��'�}�I��$��G�NlU�����6�]u��'�$8��ƙ�9�>�u %��p4��40Af�1�.k���'��S_Lƚ���x�zGN�j�3��`�'e`ٶ�����tw媓�ھ�+G栙�2���u�"c�\�Keٵ��C��,�\WJ��XZ��'S��O4�K�-��t��l���c�^C]���"��a���rD�B�˰��eS����*J}�H�q��p�dX���%�lLM�ju�4�G$�)�4�y�$���ګ샋N��4X��I�5oZ�	�3� y��o^)�x���0�w3����ۍK}..�J!(h��T�0�ݸl��A3%p⊲BFz�P�Vv��_��Mr$f�������hB���㎰*�z��'�qW���kM�zɒ +'��a37���ca�"z�hj�����2���/���ց��-�M���g�B�J�\�|>�03�qzoh�
;_	���ߤɆ�s�%w���<R�Pn$I=��%�����I�, )E��9����Y���ex+Mu[�����>������ҀcG��L�y�T��̺ԝ5)�W�;]�	�3�ރ�&�k�֣�X_;��4�#���<�J���F]��YH��N�j��Ԯ��Vх��>u"��P�ob��GF��T���G�;�2��!_����}H�?M}���v����YLq�x����e��<�GA�
V3-'���:Zl��
8��@V�;~�&{>9�ͮ|����UQ<�!�$�� w�{��{8��k�tN<��4�v��Jŗ}IE���{�|�F�s�F��N��rl�I�l;O������=VH]_Y!B�ͅoU{;�M= ����e7:��>+�۽5���kއ�I��-%Llj\tF����6J�d�Q����ؗ> 'R��R����9YTD"�L� gK�T��y��*b5tO��-F(O�s^�����D,i����Ϭ�6=�Te�0��	f�]̂�"�@8v��w�Ͼ��a�g�Eg`wy�ì�ˢ^s#��fq�@��0'F���&BN�;O�<'T.{�!L&��N�SxI��]Y�hǳ�o؍�j��)���^���H�vP��8=�aoZ:�$�z�*t-DD�Z�	��#�}r9Y��j�vV�Ə�D\�h�
�i�^2�m��n��8QZ�\Ǭ[j,%C��D21A<x[V"�41�0 �b@�|�b��q��y�G�ځi�2W���Y�.�����~�,����(#���^�ػ��Bߛ~*ϰ�v�Ѻe7g�U�����m*H�@�������+&sl��8������'�W�Ѻt=��Z�-V|���2թ	���Q�Ǧ��̷
��H[� ��~*�����=ld��Y(����Ʋ����p��츛(�
��R"���,�K��Q�� �#4իC�Wj�Z���|7���#$K�g�l���fv�A����`�iU͕�Gd�	>l�)�}�h�j�N������1�>�X�!J4�y�nuI�� t@~�4��2C =uY�`�A�z�d_B����*2���r��J`
k��i�_��gO	3����,J�eN.�ۣ*�P�'7�fLȓ����$~�@rY���㷸�vL�����i��g��lǐ��xdyKT�,��-Z��=����j��`2�kż��#�kUŤE�}��R���d{�Ťl�69��DÏw����_�_��g{r�%�[�%�1�jd��P�7�Xϑ�"m8!��$��J�����z;�(�%��Qΐ�����NNj4"�|���t�>(�<3"m0!A�{Ӵr�u@iX���ɔYX#�r��!�:OV֜Kb8}��=S�0�V��1��¯�ƅ��-<��� #ј�*����?�R�~F�{�F)4*h������g�K���%���@�?	.���X/���(�0ٸcWe�b�?%M�FMp_��e+I>Ո��j�O].*���Qgg�kl3\�eK�y���o���R��L��ap7ڙ��^ů��Dٍ�0�;�5�CTyx6����"��b�K���9}�����BMLJv�?kL�̖�K�x�K����hC�n�X?t��ĚC>0s$�i{j6�,�Ƃ?Z�*�>6�ێw�.N���IS�V�`]+Z�YT8ZBR���""PKM��+�~�����}��?�H(0���]y&�G�B���Gd�P}��BW��b%�j��'��2�"EyE��6�T8*�I�!RA9x>m=�������Yp/)N��v���y�T"y~sS��Zy�G:9�>�qy�3�Bs�L�	Q�AQ�|�#��DG
at�'[�w���#�H0*����Cv�4�hW:&��+<�>�5SābzqV���9(��f+K���D�9�@�0c�����,���mI��dPa���*�,w缢C����*�cl]�eSъ<���0��=��m���*׆��J[E(�h���4�)[ŞQ�Ǽ����i��ş��)XQ�)=���f���ʎx���x�
�̗YUj�b�jR��-��h��c�a�O�w���̿��V꟧�@����,������Xsc"OQ("�U�"���u�{�{�����w��{A��u"�l�ZK(c��s#����o�ťL9���	�+:t:_}$sV�]�mT6zD��xк��*��<CλT.�Lߞi5��ǹ�N����p�: p%".R`e��)�r�yȣ��W�����!�g��<��TX��ބ����Xy��Wԙ��3��B8�&0��g�������0�s��)����)���
 ���b/���#V�[��.�����@^f�� �������P�d�#k@m�x��Z����S�]['t浗IP��n�0��(U� ���q)�����V�e���G*�,������𲆊�(R'�K�Җf�B�Ϭ����R�&�7����+5^
���C���@V�>J��K�{�e�d�+�$�y��x�PS�r�3@��i�c��¡��ƃ�y�n Ȝn�<ɕs&#������m� �UN�n���uш��V{�=k�lc������PZY��z�p�����/��%�	�H���YF��憇�\?�qNKo�T��!�����J����P�����I/{�'v���Rז� �Y�*1G�#���m�7�M���ƨ����aAɌ&H�[?�,����:���E�Uv�_:ÖcJۆ��Qs�B��FJ���8��΅�rN�m���9��s	h�S��?XC�m��Y��.͔D�Cl��~pS�=:���k�τ�Zk�p�yR�x@�fxB��,	xp���>gh��M�ֲ����D�"4R��:e�����gX(=��Z���NoF�ەS�_����M���Π"�&� |t ��L���`��S��5��5U�Q�kw�Hf���(�h\�^�!��?Cw�,~~c�`������ָO\��Li�6�����dYk˅�c�#��	�5K���X���%�uf�nK�����[�^��j��Wi	�Zw:h񂭘������"�����mc��]�魱>K�:n��ɘ~Qr���ߪTez
��5oH��w(��js=S�k.�0��R�]UjB��m]�AL�Q���%�i''�11%�T�Ʃ�ͨ�L1�����$�?8J�����"�MM���A ��NI �uڿ�)������],�U�1��E�}(��0�ִ���U Z����.SSE"�^�,*�;�f�a䇓�X���������h[I�)-$�	:�� �ky�{�hj��w�u8	�ێ�Dp���ԉ�b3�����v%�e��ƭ��B=q�,�a,,='ΝJo�=[ ��.�q�����W�$�x#�EY�!��1����↿Q#׵��0�����*F���j����8;��TO�.h�*0�#Ky%װ>}�DJq�aaa�*���e������mB��-+�NB劎���n�����{�8��<�$��frs���e(OT�?���%j��`4��Mv�q���?�#|H؉2I:��x������8o� "HG�{���ð�Y���4�Q���8��{z��1�b�7�:��z����bP8@�'ٍ�E�R� �*]'���*]����Ū"B�i���{]0ž�;�����!
x����D�6��E�>cQ���|#E0��Z�����o�YQna*�q<�a��^͒�/�R`ݦ��4C��uG��M�*�:����\O��˯6�l�*�t�CI�1�͝���4����5���h��hw�
�����d�1���5���	M�� ��
��I�3~�*M�df1�>Ŭ7�o�pj�xk'�pvͥ�2���a�����/|���u����n��u�]���$c���r&�����?E�bL"�љ�{���PA=���u������mV�w.V��mM��R������ۀs��Zs �R�� �e��w��eTx��|���:uv��	��9���.��W���P��&U�"1��@���v�g�6�$#��e~1��|q4(�Mq:\!���JXf<=�i�/p�eq�ߝ5O/h�	����w���z�����[���@�.�6�T'��Os��s�Fh0�/�iն}Ωqf9���ļk����aeb��z�=>c�D��,]��2]te�sy7�(r�9��`uY�&�
�e���³���S�Ţw+MFv3�VM�+��-O���=aAb�`� %�$����5GK-c#N�SD`:!�{#78�qE ۓ�2�;��=]fnYJ	
.��+���O��N��(�]���������x���ފ��9x�@_-�ɐ�a�4o+؍-&Nv��&F��B�^�7�	��w �g?±sح��"e�?^�I��%{IV-�7>C�*˯��ǭr>����x�,�Y����ե!1U\k�����.[�M����w���m
R�\GR#�
+%][X����mx:K�A���mpto?���pn�pRt�|;��R��o��x��ڰ�u٭[��g��- ^�P�Q��~H骨�j������4B�`/t��˅/ޙg����S��v$�}N"�V�DZ2ov24�ɣ���ҷ&q-���A�|��P���J�Ke����g�R�538����n��)�Y���@��#�v�i����C��jOGeS�"����T�'
�ч�ƪ)5� T�c�f{����E�t��vO�a��͜Gw�Z�mF��3{ d��;��%?j�_�
�[6�'���N�$�T�ؖ��ײ�L���E���D$�訵�^Ʋ���l��3ʧ]�2������#��sM���9�ݽ�6	�b�}��D��8��<�m椃���{&~�:�ONgrZƽ���`�<sZ��
 �׵ ��=�c���0_=�=߀^_廥��ј���{� �Wh�����r�`CeTbgXĝ��#����G����%
F�t|ڵ�M$�T�M�à�(nm!��ߨC�!>U[��L	~f|�e�N�B?��0Y۹���f�)3��W7���`�C$ƭ���"�(��a�֎�a�����%��X�i�3�9l�.N4L��
v��v�����@buH��z�������a�L���̲��4@9�g�����M!����R�Ew�\*(����B���7��5K��3��&��(D��sVz͸��'6���.Y���O{$Z�Ŧ�OR��x/��BuNA���f�Wt���$P�x��o�.�;,�-��*\����,�]��
��iq�9hk������S���܁���q�Q��f�U	R�!R��7q�	�u�g��Ш��\����_/��S<��绤�	�c���O!��	bȡ/�+����@��%!�ㅤ_Z�tW�[)
5/s�����O�ޑ�^Ja�/�|�k��C����R�-�7��j�����֌�3���OhAp�����5Fs˻zU�.`��ܽJ>����������B%��(!��Pz�\U�����g�+6��]�5�H�b����Ɣ�ˌ��m�M����ef�0-=R��}Ď�'�H=� �:9��̃�>�C�9�I��d��1(c@M$�� f'�1T�t�$3��Hΰw��iķ��Q�n�^�.��Xެ7~5���ZC����47��� jbsjH���}T�
��%ˬ��A�O'������9g��>T���.(��>pG���h]����F3J�z�)qf��Ιx�'!�t��+� L�P��8�(h��K-3Uq�c��4)��f1�2"ZU��d���|ٽ��0p�ץtv�����{7�қ+�ܸ�-!*b��Unb����ԏ��V�'x�����==aEQ�i�;��\����4x%N��"K38$�?h�\�,�����������Ã�ʏR�N|�L~�Vs��ak��Q�P�0]������R��� G��������ͼk���W]T�7e �i�Ӯ�ڱ^ ̆���/�&�g��N;�F�Y�ꑂ�wҍ�P/y����7U�|����Ӓ�:�$���w�ַ���o�!I��X�pgx�Ri;`�8���9���\�|SN�
����gg�>8���%�F��{���Yw�)�|v* ���|
�U�^��ʻ��E��*�W�'��J�<���q!�I"o�֜���E��<�1�*�T�E,�|�w�a��%�b�M%>���(C	����60",��֚6	ְ���2M��e��1/����JZ�=.."M�4|�|�nWZS
e+�J%׺�k�<DYc;���C2K.��ݱ���t�5�	_=�n@^�A�13�\}��-䩃 8=2�a퉣R:�֓���>��C�Ь.ڌ@��Vl�_��Ώ���s�����"�W�qB*7(�$���[)E�[ۖ�V�K'��#�2P���9Omx���J��UЖ������7���LC�8
�x��)lJ��:���r���=*.�	^�iL��}R��Y���J*�4��%*� p�:>�P�(��@	j�U� 90��b!=q?q�@�ܐPS��	y��zu��G1����,Q�\���Fo�2RKƽ2���	���̐�Y�=��\ 
wh�l�jy�hc�0��;5!�kz�Ս 0}��K�q�n��B�Y*?5ʠ<E�83�����$xӇ�jxKs(~ܾv_�9�[�bY-e����p�ؙ���Y�(���?>}(�,�t���ɝ(^8�K�4M����Z�-S?�i����8�[;����e[�|~A&I �"C�]�Oمh�CA^�W��H�rG Z+R�!AiJ魢�12yK�@�	��JpRې�)%�,Sd�����U��Ͷ|�m�'mڶ�z��^�l��^� T8��&҂n����� ��&��TM�����((7�E�ŤǱ�Zp3T�⵳���S��d�b���E��C�;�`1�`��\^��`uɟG�H��ؗ�-y#Ӏ�A5,�f�*d��xhj�qwp���w[��8�����#T�d6�g]2�X��'	a��f�a��^)���$ЩA�ѓ���V���`�}%Iz{D���Cc�,.O��o�8l<�>�"(k��ۓL�'����M���Z^�.0=�<O��n�Ƽ"��I����l��&G��#8�(��[���g�����ej��kv���w���C���T>Oh�lȊ(F�<����u��x3N���$)�����N^��GWH8x���bxDJ�1PbRZzY�����AM�|S���9�C{E\�'��B����i��!2ĝ"��,/��4���W�X!^S�K��kb8+�',1��b�3�Gv?+�}�q����U�4��gH.@i�,��$}�k�|R����k�戂�阜1�f/ ����j��P�	_�^��W�_�i�^�e�^��jO������<$������b�vȴa��Hі����PZ�������I�H�z�V���`�($?~46d@��f;h�]\X+����a+���T�i��Z�'}�G�2�n����: H;���r��� �7[q���4Cy8!'��3�wE�-�]д�V3�!��>�'�rwZ�idwڼ��}��P"`�T.F�q��j�R��ԑ<C�g�3�<���ZS�q��y-:�!l��h�h��خ"C�GCAYӖ�$N*ֹ�Z���V#f�c�N��-/�*��k^�zY电cqĊ������ZG�>���Wj�X9z	�3R���\� �$I��$>6,f�K���v�C">04�ZB���W-�ƽ�7pT�Gq���Y½�JM��Lm�g[��#|-|�
��L{#c>�� ���/��Rt ��q�C)��Xh����<q��EgR��Y�컎�VV1�axg?(n���^d�AH��{�|�噩�jd��*�>F��b�ʅ�$�e3�\���dQ�Q�>���7�n�\�B����CA��C�����i���q�l��(�%&���?��U�;"���3[
�V�mW�XD�RK�{��}cԈ%���ѷ
-�W�%�F�$��p�`�>�ξD-�r{(䞤Pp��?"�9�8v�'����\�݃lt5����i�vH�Y���m���L������1�׿ʗR)�s1��[F]z���X>�T�j�'�7����bF �sF�UC�$O���/��T'�D7�L��ѕo�l����+VǃY��Ѷ��1��Zѫ�-\RG�?fpJW#�EO�}H40�j��L��?�ݲ��H�LZ�Yl�+�*�͕�:ј���mj��>�v ��g������Aw.A�ō�]p�.���a��/��E�2�����ܖ��[��S�e%qؐ#U
jOl߬��4��P�R�;���[�S��]WiE�����\T��ր���P���	�\�W�]xO��ʛ|C� �	ӱ��``�q�E)/ܺ�# �+���Bޞ�֞A�)�I�B�o�������^ƀȩq��;�	�lԭ��#���x��|[~J�a�{�8�N�f���pE��r#�d�ӊP����>�L	�����þ��	�Z�yi���}������O�䲙�a���Ҽ�y�GL�2b�&5�9>��.)Ԍ�ptR��Sw��9���b�1�ۢY�I��??�e�{���5�JL���C<2�'��B�����cO��c�7�W���%�D����q@+jכqa��c>P�^EЈ�!���I��%�R'C�iy��eB� t��C���ؙ8*�������i���23Wn$����;I	"��}F$n؃�b�K����9��@�`㍕$ݜʣ�i���f��T�@��k�3�G���=Q@kec�+!v4wQ��B�^��fG�M����8��<���f�ƴ��t=����~�Qg#��˒1����5�EP�? �@���Δ�KL��b��c��4C��g���O�{X�}9 �<0[�[�aX��S�&�s���Q<|Z(�R�b��-��(��In_l�8��p���S�Z��8;��N,]㠤��m;�}ȀY�d8�i܇���s�S��r��m�F��ݥ'A�,�~� ���l!Z�h��Ԛу�Ėp5��4��T�4-�#��SN<m���\io���+J�T�U���X���ʽ��O ��x��w���/�)S\Se�Mx�确4�}�'���8�:~#�ԇ���z�"��+��S�W	��^F#:�+��R��]kVǹ������o����Ϫ�F���2�VS�W��[�Ut��w?����WЄ�8���/�z�/@r���OQ���g�9�S�� gKX���q#��:+�1qM�x�đ{�#`"*ܣ�k�-_z�����{����L&`�Am�~؟mU�gx^N��~[m�%21���< �(�Y̜v�Bb�1_�Q�e���u����<�wf��_B�!�TL��Sv��T!R>�DR׮�LG�!��@�|M5�+E�&r����Ƃa�P#ޏ�1T�����^|g�
�3A�V��V��IX�y�1��Vz.P�.ٖ�\%�k@)t|<¬~��3s|�ͥ~*.��l���*u�nȿ�`�l�^t�J�I�CD��<s���	+_�m��e�f�w��:�V�6��3@��R��7���0�'G�8�Ӳ�m_��[A{}�������e�ty#;�T��j�&,��<�����N��H�S�T��;D҇��'�8$6P��G��٤�k��N�quظ��Ô�����k!h(�R��o��pVR���qp�i�,�+�|�y��uKh�Oc[�;N<�X�
�-\_���b6�p���پ[�K7U�k��ݧ�)�l�۝%���iDg��J�}[$��G�A<��S��1�/��OeF�����Ֆ�9���폆L��~p7�1!��{<+-��إ"��rK��I���9E����X����}?��f\�l�2l�J�|o�!im}K��A�ɺ�̤f��k�0��힁$�z��ܝ���o�W����U�\�~��W��= 1M���k\�8����TNgy���>pqP�)�;~�0E_5Og�=��+�n��$��]�{�
<�(G�6	 �0?�뗵b�B�K��!r�O��O�X��7Qя�?��&5OkCm�����b�!�Ɠ^=_Z�Pwq�rs��C���Qme y?�Ĩپ�����:t*�`�1Z�� R]�x,�m��XU5Q`�~���֥��S_�e�>_blD�2H�
�c]
v�O��-;G�~ #��r�;�߈m����h�?A*d���z��RÆ����{-��w�q��J׫�<��c�75�F F���M�^����K��.�Wq�*AT9po�L�5�ҌS<�&~yu�L����G��K<$b��9�R�Ef�V��֤[G�PƌZ��eI��L��,�5��Nӏ�+���?SR�Zތ F|������R�Q&4�Պe��F��7(
ے�~f���.�-�Y��1�J����?+���Ӷ!��
J�mfo�&�S�ib		�5)2�C?�[���nL,�<��#V����c�np�������O��P��Ҽz+�X��{����`��,�"U�m���K8���gJL5� �g��&����f��׶�2��e��X���-m"K�F�j:JonH}&[(��}j��BΤm鷒��_^�ը�a��3��~����tX�乊���Gȱc��6������1��#3�Q��<��p�dnNRM��S������9L���/�H�����P���o�ѭrDSe��Y.�O����M�R]S�)����L��1�l!���}$��敖^O/,@��5��j ��ԻC�)�����z�|�0�Y�/-��ᥬ1�T�>�V~���@�OX�u�,����9���9���N�>~W�N�i8d���:ŮI)�~���Γe}#}��_���*��
٨̑�a�H��c��$R��4f
U�%���ɣ��Hd�j�۠��mwJS��;��<�?���y���UP�����	�z�c��M�y��H׊%2��_A��H����-�LW�N�-C��gzw��[R������(z�}���u��	2�K:	溡3�ah=j���TU46�d�c�O��٨�����>���;����ʣo{l�o��P�5\'l�4z��31�� z��	�0�(�2P��'��F��CZ��
� E�����>P����Ϝ��Ɖx�Fj�y0��6�`4�A��� �,����8�Y��E/��ޮ�\3������%�tP/WD����G�� ���5�MV�\EVkt�=]������O��%�l7�������ÆJV�'��f�P�HX௞Zʥ%T;��E�������������X6SR��ʑ-��3R�l!���1�mF�F^BS�Z��=B M@�e �B6�3��q$���� *���R����y�LC�dc�z�m7����������U�2�~���I�q3l �&��AA�����o<	�,�7�mzLMY�&y����w����X���	��v�d�H��� D(�?=������}��e6�1j\��NtU��֠����4�ՙ��'�	�IqK��
�<�M� d`T�"��9^:is����:��D�+5G�|1���� ��VKlt.g��#�ʼH��>V��oRΎ��rw��g������w,:pn֑��Ǔ3�����\m��̓j+��Q8�Ճ�������<�R�?5$�Sx���x�*fJ��Ȩy��'\���Qa۰/��pj�@fz~�M��%����p3�5���l��7�.��Q��0�g��H�
C�O;34�o-qF|m��½��ð������X ߣ:?�[���56��ާ��ꄂ���!��(�rި�������.݅V��n�J�T����En!��irX�9�ÞC� �D�6l����3�L [�P�����}�ׇe�*FM�1m�6�W����yxK`��v,��،��j�#~C�1��S���~:��`�~�H�_������J�\���YC�'�u�K��1�lq�L�~ .�6�vR�tU�ϰ�+\x=��F�?f��9@��������i_,V��қ��J���&��f«�n���tU�=���dn�)��l�$7h�� _�Z���<�i�9��%͈�ǀ��tב�c=�GrD6 ��hTJ�BlMP�Wv�˃~������a����ы��x1�/��@�9�Jlo�Im\�h�L�)��VH�5���ok�UO��v�6"��������G���@4a��U-���:4}��G��c�n�����q=���7�x2�y]�:��H��w�#�r����N�l	�q���h�����׷h�^l1��	.���`�b<���g�%��м��=���2������G?�uwA��]!\	Fg�)��o[sF�:��sL�(D�e3c�^)0�4�?g�8�����
7���G�&�m���D���U�����Q���O^֫��fD��W�}�F�1&�>U��:��nD]r������s'ż!��S����������
=����i�� ��)��*�my</�7��K~B��d��5d��N?tp�-)jU�� R�!:z�Q�-j�z��rP M������� R�2Gڇ

t�P�rɸ84�	�o�:7x+j����eK�7���K��V���P"�{���'1�1?Y?S;'�|nH�=�}��A��|v�@��ٚ�(���`�#�Ē��~%7��)��i�}�L!�5L���ӄ�8��f�ʑ(5˨5��W��� �V���q!�Ԅ������Y��Źϲ-����V�����5�T�w:�e�$P�I��(�m�x%c�o���쿐��6m�Y"Ygɥ�~vn�O'�1j�����y_�p����T�d�X�j�J�6�NV�k���.�Jt��A�}I�=<�������b3��m^&J��BQi��Ǣg��♹ά[�� ��UUR��Vg�Mg����Zn2���'chI�#5�Q��C��(
w�{0�L�~$�i��'�p!*�o�?��Y�7�F^��Ƅ�"��g�:$�&qv@�L ��ym�G�����g�7�������9��H���e]���[H�����3�WM;Y��!r�pп�+�}
F�B��V��@lXM��D=M�}V툉���+3�y�>������y|�3���8l��
Vs�1Y�� �K��ۆ8����Pl6�zB��S-�3�h�>��0D@M|9�qR�����g8h>d��pR�^?��~?��˦�je��V�!�9�)z���ٳL%��9Bf�.����
��,yUFs�y�B�1JRZeG@�9Ў�H]a�����L�x��dH�
cqRCw�u�T�X�c]^(
�]v�N
��Ǩyf|.x�U�D�p��Y�̫�&�A'�>�E��H�|���Y�1��}���k�0=Qc�8����/*��L��"3��c'�k�ѱ�HL�8,��7���vN��i��2������E^��aWH�=֏� ��ݡ0@j5��r1%}�0UY���k?�e&3�ƽd���~�^���-��X(�s��,��.B�i:��,�Wq�}���'@�p@̱��'A=@^�XE-��깔� m/"ܮ}����^f]ˠV��i��zK�g��U;c	3z�(�Dw��S"�E%7��^��d��VJ��9��39�.��P����Y�
W�fx�#<]M��V��3	R.�M����B[ƞq�}�EC:�5����d�C<���T˫ �����r����j�]�s�Ur����U1F�B�j(V�`1�1�l+�͹��j�mt��D
�V�Ue��ۃDc�p�c���b�4�re�h���h�0x��SK��*g0�����D�?Ϡ�bh��CL�������M 9��o!��'�.B�Gp� ?��c�v1���#B����u}C��+�����o��v��U�� \�v��~�����a�9��f���z�gk�<��K��!n�4F�k�ԬJ�x�|5�Nyq�0�iQ�kݶ�X��w�M_�Q�M����u����/�ǩ��&��?��A ׯ5IZy�ޖ���6�r�O�'��q��rm�]�'v��� �1���uJ�1�	G�[��m�n�Z�� ;�._ȂH��N�f��a��N�z}�����3���j���5MF.M�ݔwR)���Lĝ��}�g#e�n)5�e��v��eW�X�C�U�k�*?�le�Q�쵽�V餁3~O�A+0d�}o6Ӹ%�oZ�7���R��Ӧ"��C�#hti;ÍA��/!ThX�+���4�n�럵1M�e�KG�(��B�NR�f�����H��ޤ�6r��u��$���g�jX,P���K��F���s<OY���Ґ�H"�n=m�K�D`��:e���+�&���1WtdU��c&�H����U�r������gl���>�V��$�;�?%DY̻�s3��sLn��&`��7\<�1����N��JZ��V����$i�治�B�'��^2���Z�c���"�Um7���HF:I������i�� s�:���c�]�W"<n��@��k.rj�q�pC�������Jl*�Q	���u6l]����S�,&��@�y�(x�� �D�(/����f�	���ܷ{�X��ț��`�QEϠ��i6�}�ds>�,�,`�@��<�M��^�p%!)3*8���GF��4j�N��5�m���Or�:M��kl�)k�A���w�?�����*L����8({2=�����[0���]$��5���P)�wRpm%��V��r��]y�Q�cZ�[�t�*7�aH;���4k��U��s;􏽉��lkc�WY�f��V��/�L��#�)mP����-����_��̦8������^����b~�P.L����Aݚ�+շ^�.���#��NMD�ް=-�,�l�wfe�3��;����/!R���0t?J����%�*a�y]��
�mp�i�\#d�\)"l�!�A��4��M�w�v�g
e�@�E~�N����ۑvZ�*��"�9��Ci���6�=�8+;p��E��G.3�p�ϓ�e뤉����b1�56�}i��@�����e9*��j?_�3�E�m�L�����|�2��IP(*L��R�u�� �V����� ~��Æ��45%@�=w��S�BN>=��3�mp�� ���ُj��R��=��ٴ��v輵cW,g�����zy��!��`�T�z��V k�=�o<u���o�e	{&�a�qy�\�ui�b]2�6��C[b)��{ݠ����
&@k�F�x)Z��钡8��ǡ34 ��5h��ϭ�	��R!	RW�?1>��+6@q��c��jwL�<��`���̈́NA� =�����[]� �6�S2�4t�`"���5�`�;t6����ѝ���'#��G>�ښ�78-Cv��4A�8"H����)YRI�= �#�Z�W�{��GH�&�����˵T̊�n���nr��8"��	I�1�ʜ�4u��Pn
�n��%����n!t	�Kh�m-ڮ�~�;�V�sq��
�owVn�2X�4��瞧d��z�� ����"i�2V5bŽ֐e�H��@�ؚ�LW�2=}��.�1"D�TE����-_��fm<��L+�u0���$��ybp��
F�cM���[0�GV#�Q8@;Ѽ
r���	2 X7n�r}p��a�?��E���=Nv��`���[	JE��s��57���r�ӦJ�?��wۼh�� F�!�K�W�bpq�b\�����ԯ]�ѩ6���A;l�^��[�z����D:+�뙝Tx��G�[$}eI~"�M(��f[��y�UY�N�Ui9�Hwn�%U��;'�d�B�D�U��	�i�"@-��ƴ��Ӯ��p�����日b���i ����H��U�F�y!�)��=�q�vS�j)��?��W�6�=z�/�n&Lf��.}�?��$u_I��/�uQӸ�kk��_@��� ��������Pj$����S�m���u%=~R��3Sd��#��'=������<'I��|a�	���U�5�:�q3�E�uL)pǔ���V�:f��	��Ӷq�n�>E���1�=�k8f��[�����8�LOG�ACY*M���T)M]v� 4���N]4f��j��/�3ܚ��y��b2����A��JV7je!Fv�@�U�#K�%Ne���d�攨)�Q?�e5�� ��2���W�yve-}��O�!���K0���7���H�N���OҼQ��ʕ�i�@9Q�提Kb�)C?r�������1Ц]�H�|q ��Vם#(ܣ�i螄�[�������8�!˻R[�,� �v@c\i�ߒ��f��]N���{��W�f�."��ލHT���"3��]��W �H[����)[O#�"����ը�tui��G�kgE��;a���Fr�
	Ә�	*>��94?����d��Μ ّ񴚂(C�HT���9+��ƹ	mѢI�=&������H����@E��FVA��gl6�~�mI��?���3��i� �t��V��������!'{�+Hj��Z�FD�0Vx���/Z��5/�a��iaq�`�$��Qҥ�Zɚ�y�6Y ob��?��oLk1�S����c��꿚�r�[˟� �㵙2��'�e���h�GHh��K`����^� ���.����0���^�	�}�D����j�����U�Yd��x�s9������}��k�B�25$h���|�\�U�纤��FD���d�H�a|59�3���5��Xbf���s�0x�Ҥji�Ԧy�&m_�TT~���q��ڽ�!��H�o�g����&��Pa�v���������ӫq~�Elu��O���-�mi��_�J���@�"Y��_?�5{=Jr�`�,.5N�{�ܨoWн��q�vQ0 @L�wJ��Gp޾)G~e��k�$U��V���i�G#����8(��Sg���;���E�����ԹU���8Λ�ּyVM6���X%k������G���a��N�L5'�{��`A;��UO��$q��H�z��g��:TT�2�����)Ȇ��r1bO*�L�my@��+�q�:Eh�a����,|�b'o��� ��k���zb��5�6إ7c�[���xe�[{��x��0�9!V	���ȶ�:K�
�Z���� �7Z1_}B�Q����S���VO�qp�2���]�;��e�:����jI6hs ��P]��d���0o��#v'*����<o ��LV��䫦�o%�hu����4;��i?�3k=���@+���ʐފ�u"O�/&D{��t�6�H�BL2�}@�$ƪӿ�y�ޫ���:��ѐ_�^=�pқ�*�o��H���R܅ܲ!�Pg��Ҝ��{;��l�\u�����"�e�|�JSi�P],CԚ�P�n�2x��Ȝ|�����\^�:R���a��q��	��%x��Ն���b�BWk���F��D	rڀeu<�lHSמAϘ���l¾���Ȳ2�K0�����/�6^{|F=p9f�1��A�M��wR:w�C㾸Z.�B��Feg��������7a$J���p�;�7k���z�l$�S@,�5֠Q�ӳp�t����������h��$暢�>�+an�#4�y�QvH̆�W�Fn�.`3��I�����㍭�޷S�����L�$&rO����ȧ�I`R�|O=�	���!�<����ĸ�fպ@ͩ|�IR'�W`�ޝe�9 ��ZP��틇!�m�g���y-�!���oc0=�Ȣ(>���e�kŧ��`�.'n�� �����=#3�>�i�@�e*�[�L��	��(�1�n��F@U�vD~��h���8%�5
ҍ%�̖�Uo@.����� ���?�C���Q@D㟺�
�0�#��r���5��祜�!�FMv*S�WK�v��&Bu�6�eS�@�,^Otj3�^yjUX�V
FM;t���\�M�Frh��w$��e�Q��G:$]�7~3�c'}����,�~��v*���C�i#�����a@l`���0 �#��YOQշ�w"{�D���4m!&�����i쑰�1c"�kCk��~��%���+�̥�m���I�tVY�#��R,|ͻ�K�������q�y+P��r���q"��Vzg�ko�x�j�Q\�]#��M�I��RPt���7��i��$�3����b���^-����B�y��S�eI>*�_���5p?��Ϧw[�"i�'���g�Is��:%�֫r�2#��IgMG�����8�xdq�}����Y�7W��f�q�0M�^��٬И9�7�oB�s{b�ʓ>��Aym�0�B��w����2�[FP���rpjY����Pp�	�[����t�rb;Ek�F�M����U�v|���Z� 5��VƢ�����K=���?վl��Y=[���l(�f��'��b�IwE{p:�X��1'BxɃӺ#=P����[]t7�0Q�0��O^�����^,��:s���3A�P2�2������RoY���
87�g�H�2��|C:�4!X�jPO~؆�D�R�2[9� l�oZ���<�Z3����{����K�`��^�EG1�<QjT-K^V�|��Kѿt���}(�gK��~4�-�����W�&�VrIG�U;�O#�A��WE��;���|���p@�.������,���x�zVj�f��q�6H0���`�>��2��+D��HDs�l�� �{�B�~|���q�
�������=���]B5���î���;������IƑ3���[}	V�W,�$�����sL�3��ƲM5�=�[�/���L	J�@�@�_�r�E�\�Qk�o��y7�l�M�a��k��+�r��
}�DOs�Gd��^���9J����n
����xQ�� O��@�OF�	��0Bqi��	Q`?d>�frQ\�q��/6�J�2Or�g��r=� �l,YG��o0��f�KC�^V�7*���޹�I|(�y�D��~G���A�0�6J��'宠x��yG�b�qU�`��Y������o��2v�H|���v���}�t��~?���F6�:]^I)�ℷU��J�i�c�,�N���o�4�a�8b�iH�y�eǉ�Ѿ�j��^�jk�&y��R�2�V�|X�]W�2�4�C�K�G�@�֘���2&�)SO��j�5/L��)%���i�0	�� ����WDý^��^�8p�Cߕ^fS��·1�W6�Q�N�n��;r�\'�17H����T3Co�[x�3=-� 2#�@%��D�>�@k�@�N�)+F�-Pꋾ2�7�y�������m�7h����_�P�2y�O��g�\T�; ��M�-��Q�`�]p��'.}ㄣk��&��2^l�-H�T4>�!�U�墉� J#���O%p ��ԴI34�����m���l�	�O�i~��S������2��P���+�d2���g������kY�ڱ�Ѥ;k��C���ֳ�YAB����0\	�O]?�L�[˼46���cH~��"@33�ቁ�{�QkuE��!��`�w��[Xr��o:��o�����v���Zð�j�`��!�&	��lCd��3��p���_ǧWV~�M��70�qO�[��Z�*����߄8�2�$~�ƕ�
�z
���)�˹{"�"&?K�؁y�.���e��6$�g�鄧X�Ֆ����
�wRHL�m�����m��5�3����4%
��6�����u�*����Ǳ6�����\�T����6CA��.ي�����0|�*�5&e�VG'	�E�f}�,����݆�!h[�Bܨ���.�Z���@�q��k�-[�~1�v�]�f	�M��0��.a�$���\�]JO����f�_��؜:�c�Q:=�U`2(ʍ~$7�F�+EVz��J�CV��ة�,jʳ'���S�����?L=m(�R}�6�o�ٰuҠ����2S/��Դ��9��U�IH����t����W���]Y�ӌ%y���M�W'�bJ.+d����+�S��X?��ee}�.��u.���#�L!.-�2���<�� Yސ�nzמ�h�sM�Ne`���+ �uh4���S�ڹh*�H�_�_?�@2Kb�Q�c�뭴f�(x�2��������Pgq؋Qo������2�}���g�\N#�m`.��_��3gu�L��1�aò^�)�e��S�\�O��R?�Xm^]e�bs�/@�������ᖚ�އ����?]\�O��7��ظ��7u�rM�H,��Y2&#Z'f�KUO�b�nN�_8M5�CM0���k�Ejւ�K��v�M�!��V/.�Kp���|�,�i���m|R��~k�t<�o��^RG<�Cݮ�y.�����@�bّe�^�y[Q�MK�D��7}@��!�1���ā�E��iY��C����("'G.�cͅx��J��P��HY*�?n!6����v(�K��H���7Cw�	�J*�[�QuUUAݛ��|}YGľM�,-l)�-�$'Nу�i��18GO�44��/��w�+�K�����ow�HF{�#+N��F����n<���hj����!���~O ��Z��_�%��]�{9\k�� �ϢS��t=8�0%k]��|��8�DC�[�i�\fr"J<�PS�w��o"��;�k$SB�����cs F)�)��t��ձf�gJye�,������fF�sL�8�0����������:g�$�������d�M�A�O�0�G����k��o'l�����%vM�GU�{�7W���y!�c���P���B��&����cVu��;3#��a�����k!O�i����8j����4�ng�>}��Ŏ�S�n��)?}�I���ai�m��Aݪ�n89]���܂�Os1�E�ڈLw%� �+v����N�@�@�6�.L&��G<n�-�} ��^�l�5��7SS�g�$S�X!��"Kn�9Ƶ(Jjd�t��J:�/n�B[V�����a*r��\�-���p<�_2���.�Ӳo���GO*K~W��~��  U��U4%�Y+Q"`�����Z�s�ERm,��i��g��XQ��SmE�Xh��A�ճv��ǖ���cL��h!}	��!�^[�߈0{e���h���H(��qj�sςKKf�2��PE�4�F�L�g���;-Z��ۧcy��A�0��y``3Ss)�9�Ʌ曔Y:�ҥ���fP~�6�WY bj�i�I �E� +9�7-���N�z$�L�H`/I���t���=k���HJ����IPd�
f�_N��4_��\8:�^wυ�������5�H�v�iZ�`�$���s�д���W�pv�*�:�p(����5��X��y6�NÒ�h�w�8� ,�@H�}���P�8]TҬ�3���&�.l�8��3O2	P;vֆp
L��w�@W5MŁy�I3�G�U�kF����FX7�Q�.�-�!�1A#��Oe(dp�6���|/�C��R��w�Ӌ�E���Rf���Gw����=1�oyr��#P�%Ȝ�QT�h���L�.r�O`�u��x+w��xP�?5j����xŧ%-��̃q@O�8_K��SR�µ�"������0K:-Wy�&]���ϯޝW}�hX/߭�����`�՘�+6�j��&�Z�V�:���~�Ξ6�s�L����l��SV���V�Y�*����v½*��rG�ue�4u�A��gA�8�4�h�B���?ho6�G�}�]P��f;]�
`��w�J�-��l���M�Z"s�v���&C�Vв��h�u�0�g�=�i�<��A���L �#� IE܎$,Ng�B���ƾ�u��0�	j��=�G�L�
�Y�S��e�J2����7��|�gN�kS�@�]��NF��s����ӿ����0�\i���фn��Ԃ�8��uF_�k��P.+:E��@�T�Kڋz��S44�=�-X=݋��[�܁K��!�;ѫ	`8��Hf�o�Jy&{�!��X  ��A<��$U`�-=Y����(����${����(Ṣ��*kOB�m�뎒S����;�Q�7soئ � �AB������c�5�Ճ�0�+�<
��~���Q�ֆ��������z�Z)��C)ݬ�z�������"c��L� �A$��$�f����d�c?"H޾񐨡k&��oY�y�>P�f��x�X+����F`�SL��[[ �$T��/r���d�~+����w�z�M}�H��B���ղ��g�KR^��s�Mlw@�MpO��=�7N�Z{�ﵷ�c8�pr@GbD.'ۢEj�M�[/�f�jAW���J���R#{��8�72�C�A�xr'֊�!��A5�dF�"��9�|�Wb��Ҏ���w���8��np���y�'R��ҽh���Ě�H��}���q��%L}ni c���D�od�)�x�t�=�3��w���:�fDsj"
A�ףı�(4�h�N�8�!6n��ڌ7�!�f{�6���|���J.��mٗQ'xX'ҙ@�)�ú��ǀe0�_�"�kb��\��w�L������uP����+>�%D#}F��5�5ʡ�J"��z ��r}֯
|��Y(qS����o��ѢN?��£1��xO��4�GQ~S�3�q'Ml��!e���T<ۍ�n�x3G�Qw-3L�������\}��TX���1���k�q8�O-�H�-��
�mV(���H�-�o��������Br��6��M�3哃WN��݉�/Ap�s��L�+BANc������̰O��P)R��QW�=������Y�Su��[��u�rRH�8yy��p?��b�Ί���dؠ���A�6n�^�f♮6�p	y-��K���ڏֿ� ��P���ǧJ�I$I[��ϺMI(#x��q��p��ʿ�C�L�|"{��kbC��p��hL�ؽq��� @��EB��bK��B�M�)��E0_኉�.�Ӣ�`d��g�a������d3Mӛ��O�P��ݝe��̩�k��+��/?8��nd�k���H3	�Ѽ�%�{�dw�`�ϱ��S���|&34s� b�B�!
��eI�����B�Փ��A4�2FR���÷��:�&�!5u�=sn��(LYK���H���K}0g�[V���g�S��/	-.��m�#������M�P��¾�O;ݬ�la\S9��5�*�pT�@��[�P��h�<����H��Ŷ:st`,��:��*;7�R���L;o�F�j'�(u��4i�hƭ���-��i=Y*���	A|�dɉU}3s2eQd�Û$��Y����F���}�I#�>b�)(���|) l�Y�M�O#MV�d)�0F����0
Zu�0q=I�}m�m2�ψ#��aM����a�m[��$��H]g:�(	,��(���ᱴ(�&�y'��2�I��yEHR�B�'W�q�`�"��d���lt��{eϜ_~Ϧzs�� �Æ��Ok�Rh�.8��wSo���-�R�Rn�"$�ވF���6'��"x��1y՟�f9�h"����	5�!X���g�V�����W���"�Ю�5�:	�2eyzRz�!�&�����ޓm�U�ǥb� @հ����v������H�x*�Y���)r�n���G���7�'�zd��1�s�V0��x�)b�e�)�vO�k���TC�:���/B���	폧+�p0/$ �i���%��E� Q�{��J07?�݄���ݮw1�DH�f#b$&��� k��=�I/8�^R�9�[���u�nbe�t%A9y�NB_��%y#錃��o�GS�}�
^*uq����:�T�N��l'�)b�p�_d���˗](��x�q��j�ͱK��B��7=J�4l×[���f�O��[M�#ٞ����Mu�m�����b�DoM2�Cty���	|��z�Z11ʗc��E֥O�5M&��U?<��L^��L-�l�;Ծu����v�v�ʚ�k�9�x�煎�0>Y����4b�Fh9�bU:i I���|W ��:y^�q��E��<�����njY�}l�y�X�R��,�|m�%����3�{,F��7<�Z���S�����n�5d1�Cf�O:\�󋖉�
υ|^�3�:þ�̗��ۖ�l2c���wq�����ԫu����r�'۝ԇ|.����-���p�җ��(ppʢ$�C�q�lFG������P踷�똚��x ا�Y�r�i�m��x�0�>�� :$g���M����r��� #bp{ф���d\yU��H�r+����+� T��8�(Uv�����H/����"���hnJӕ(@"�A���8	�lH�8D��p�{Yy�Zz v9^�➺���HZ���I���d�C��v���2U��;�� E�~���R7�&�4Ů1_.`�s�D�5H���ZtM�#����T;Iꊅ0��G3H��(@Q�%�u��z ,A�a�r��/�Jі�gb�����YQ�����)!L����:ա�O��o.L4�w��	y��?���Ƒ�L'��	�o�z|��&m�D��`��P��@]�v}�>���m�M6��t3����� �I�'�L�H�Z�vA��9Qw]`r�z�SIױbٜ���/<?�#��Sc�L��y�[�^W�d��G
�պ�BjL��l���)����L�&h�������ŏ�G�|�}����AN��;�H_LeY̯{\ҩ�"�|�NL|�?�c�B�t�(��
�Г��> ��S(�$�}���x��/�N���	'�:�A�qи�y���TF������x-;��y�"X?��/�
��j��Đh	]���^��eZFs�����A��F�S���ل�4"�����R�N��i��G�?m�X��ӱ)�/�a����	��ʬ	_a����h��n��E����Ѱ�#�P�b��5�����>Nޑ֖gg��T��ֽ|�LQBJ��7�a���o|�p���<���bB�M��d��F.+�����;��I97yX�`�<��::,,\�{�>��!�ΐѿ<��t�?���J�qsH�mQ���=g� }��_m�`������&��n|�L�����E�:%HU$=A��:��76{��;����L��VD�i%ZR�kY��4M��BĻN�^�֘�8�R�]��?�>�����f$�`�ʷW�7
#S՝M4Cc�9��J��"���K�@���<܇�RB9��iNW��6O������RI1TD��||��NVvc��Q)JE����f�x$ ��h	�!e�M>mHZm���Y7L�h:�����K����
�{
����q��5ARr��)W��b���	��,Ix���9�	k³g'Z�����V��迻��eedLS�QH����jx�����'�냲r������[���k�"�.�OC�qI��@�M�Fi��NƇ���,�Y�/�,�[�Ӹ>���MD��m���z�@�����`��<����~���c^{�|�C|�f� �P��2_�Cw��V
�ƺN��U(�H���#��Kl`��Ű��2+��1��񐈼� ��lmH���T�Q�@#}'W֟T�GUE�sփ$��P��akӯ�Z
>�T��풀HPp	q+%z�������Y��,����gjP5�|�f�\�w���/�﬒=Xڋۼ��?\���bY���Uخ[�ϾN��#���M)���K�E���������s.�0א�s^��2c&��Z��7&W�����X_M
Cv�\ǚ�%�c;�S�%<R:qd��ɫJ�4�U��$'P�ȕHT�1���0��>;�q�?獉���S�@'�����o�"���+�����y_�U{s$�����\3=�;�̀���	`F#�voS۞��UU�#�S�8�DL�|��ȃV�8�z��*+��#�V�ګvI4(� �=D�+��쾅�xoБ=�E����ר���c�&Cbɧd�Ɩ���B���$OY�P��i��7T����M�w"��z�ܣZ&N�7�����]h���'i��_�w;��g�ؽ�']7��P���0�>�?y���a�e!�Iz�:��L+�fa�ݰѠe��fE���~�#��9]UC�7����@��AH��M�&�X�b��l��#��dN�J�����P�	�]��A�/c��N2�Hs��t�z]�	�dӜ{���j�p�#�g!  �6�� U����F��VR��u#g���RsS�7�F0>i�y/'!E�z��Q�éв�@���k,6�Ni�Qi�M��&�3�Fw�"�n� ���#
��ޜ���g�/��@0�Rd-mP|]����rr�^w�Q3v�HYA��|x�h���o�Ef�W"8�Y�e:g�v(��-��G�p��DL�L'Br�:����76��q!�뻰YM��O0v����'\N���5xL����M�B���I �쐗���kV���|D�6��+L��oI��Y	��Ӕ`"�]�6�qK�d� d�!K6���c_��k���b�p��n���t�5��D����fXg��I��p ��B}�)�"yF��j�a���o�h�n�mۜO�����lp(�̥A>Z*g9�j��q3�՝\��D�׍���PyC��ݐ�W� D�%z����U�So�ܤ���YDM�g�i�*55N����M(0�&���s85�ۀ3����
�[٢{T�x���:[�<`��V�r���5gK�\0�[?�c]�ڬn�����
��{�����>�oU��6j��r�*��O��Yɖ1j�^F��R�FG1�bAo$/HY�<[�ȡQ���hfD�]n�����;��q��pwq"��z6�@�t,Y��fm���P����4�A�N[y�&ԩ`n�J�S��l�.Y<s?�:)\��
A�v�%�6��א���N��(�*����F2��7d�C�
�kn2z1 ���->"oa$�ǉ�YZ:�`���̩8HπU\Rr9��	c>k{ ���_n��Fn���z�?}�B��Cw��ĴAՉ5������j��W9���E>���k�կm��`9d1"h��h?d����R�T��Sq=AT���TEPu��F�WJj:yu�B��$�K�=9ʎ_g� ��;u��4��_sR(�0DI�q�y ͤgg9}t��e�Y�kL�Y23�"$c9�5�	�d���9r:�Ǥ��$�rE�c܏>�7���K�I(��u|�ҁVoa�:�9�hD�#��� ��>��L�?��$Y%D��r���CX(��Qx�?<���9x�bͮ�ת'5�@9����:�<J_��J�4t������CX���8|�Xa�� o�b��F���&����W���%��ё�@�ȅ9/���H��Yִ�(h��=�q�l�<�Y[�S�K� $qgG�sQK���)w �����"��j^"��-ƭ��c�1K�0��]�.e�ܒO2J������@�j�F��#ZW��t��?ޢ!48<_�\�_���g��B��;ݸ�1�oTo�/�ˎ:��(�G$�����a����7�w��V�ܷ�
�7�{_q�`t#DM�pLi6l�`F��`��D�u��e�;k�^W�~,ȶ}�ssK9��7��Z'�a��o�Y�&a'�)|����-	��DO�ׄfk��1���Z�q��ي� �B��bx��l�׉K��P!�d�q���۬��Q����ŗzwӱ�0Z�&��ع�����ķ��"�	Akþ�A���o�8��,^IL���9}}���d/�5̸U|Jc֞B�����P����KD$L�3b���
�<_��H�Od-��r�^��j٠��N�X�b�����s�oRy���i᎞��2�|�
I�eT@��dr���J�D9�&��U�����u!<�1�;8�u�fJMa�6�5~�%�O6�,[G�A~��fd���r,혥{��A8ՠ;��T� =�����.�٫Q%)`ma�3�\��?F�/;����Jw x�-xH�ع���N9�ǎ�L<�g(�/�S��\���cOj�L�}�ʛ���a�%���>0vh�5�+[�$V��e���ʇ����4��ʽf1�������Eƿ���/2F����n�#PS�6���\�mݫ�N��ék�l�) 2o!ᶹ���� ���#j���Mf���F(�ӊl�Q�@�s����ݑ<�@|�ַ��RC[�s?]ǠS�W:�CS5�rJY�t�͡�%͌���!�Й�X�vK�0�C�bZ�_Rt�/���tֈ�0,����?�����O�r�R���NP��C^A�r�}�BWy�&'@T�+g<������u8;7���*�(��K꽓����	J^�K����v��X�B}�˽���I����oD�g �4`�����}���=�꿼�(�c�VsM�^r�C
JX,��iʥ����4 �;��p����-#�7��s� L�Ce�iC����"��؃�  *��Iÿ$\��V��e&���&�
E��l.���o���=u *��?���I�Gz�9�ͷG~�P�i��Z�tvȗY��n\����~JK�?t�4t�څ���U}�����x�*J�IpKj�H�ڜ�
������.��������2@Ք��6�K���H��c���Y\�o�.�+*�+��Ӭ3��!յ�<R0N��C�]�jΒ�]j|����Dl����-�Љ��V %oޝ���(o��s$k�3��e̛r)%�`�W<�|AK-�*F�f?��Hi��`YT&v��m�Q0ap���Z|�ҿ[SM���o��z��tU]�HW�Ԡ^/-�pMR��A��lG��`���L"؞"�z��.$M�w}ث�������$�x�X��Z�˒�#�l4�@�KT������ ��ufe7ωYF�Qr1�Q�?�R����ζ8������<e* ���#:�kCdTwx��~e�%�:�I�#����U�ڕі�\Wݍm�%5C\�l��kLk ĺ{Qj/h���/�%�QY;��!E�9�oT��>G[�W�r��f>�%�`
Ǽ�Ev�����D'v̇ºpg��F'~���"G9����xw$:ŭ%>��E�����1���.�~��蔪b,�HWӂ�_��:�mv6vI[���EJ;����-b�4����ϵ�1��b��wt9�إbjE��Z��9����cdSng��t�F�����?�ÑeG�WƠ�ݽ�rjQ�E�چ#4�Z~�#�#�ef�ʅ��4 �'�v[����v3d3߃�a5y���s܇M�w`���_���}ׅ�5���k9����)�YMb��ϊ����(&�t��q�,%���`),r@�b(�A^wY�_	Z�6N�{\`�|�Jh�.��$�}*��ȩL`�������`��@�'= �O=�|e��Z�\��g��?���C��j~F"^�y%�c�O�Gy�ݢ8u�e�솄�!���������r0HC�[�f��|����+��Z�N(�%4+��O+[��8�gm;"��_(V���ڋp� ���ԧ�xY�B��	��	�� �e��Ȗ���n1��K�;<�n�K%3���uBɲl�OV�����+�u�u��~0�e�m�|ݡ�a��99�C&[L*w׎"VV���g�b�=�ug9����Q��r�4Y6x��l��Ŝ���S�xq�{蠎�ү߸�N�%�x�T�~$wp�uQ[�U����F��د�K�x"칺�f� ��5�u�It�M��4�챙�F��:|5���%�Υ���+m��pg,���^���d�ؑ ��kV���ܹ��=�[ ��V����苊��|"6��ﵴ�W��AhN�k��9�MfJ��LZC������*�ԣ�񙐟d'�>Ce/�L��J��H�6	�%��Do4��q�P��`���e��5�u&�#!�q)
l zrb)ʪ���{d��k[?�;���v1f�@���)=F�L5��_��B��e�W�#�1��J�Dw|���dҸ��>T~�z��5&'nnU���E�,��nzƿ��l�w�Q4(Y�
:i�ah<��:�.W�6��J�U�]�h}^$�bJ� N��ɎljwPS#g}�Fö�o��+0�Ie�[v�S�?�������#.bb��F�69?#�d�-����x��z��5A�<y�fV���U�O�y�-���e�lx��)��ܤ!����u(�Cj���nK�Pt���[ ��Νw�m{�Qչ����d��O�a�K^B��Z���bp��JCəK"����,ϱ-i�6�2�1�#��?�5� Pn."��<�	�n�,<rK�_�����zF�x�h���a�x���	��AǼ	���,��:/��,�U۴��������v�s�C��zk��D�X��ȭ��M��	�$w2��i�01	&JVh�$|Hl$A�c�N�1��~��z��O��Ӱ(�<6���y���fm"�e�� ��eE�ؕ�(	��z���zM�J����NF'�c^����z�^�jW#~��x����-O�+�!+~���<f0GK����'�8��;�9>Ga�rъ�yg������	���QG�*��R��ʹ��o{Il%����"�վn��uR1����o�T�X�}���"ɓ"i��lE`���ێ����ե(�����,xm^`�]ME�v� �ܧ��0P�Z�4����+�.��~I�Ԅ^C�� ���бm����kw���X� �d�e(��;���Ĩ,Y�xվ��U���5V�'P�o�O��X�k��Wh�ǀЖ+TUеTG.���q�Y-h�ɚJ���f�{h�[֧	5=�i���m�72@^'Wx`j��� ��Q�:�cZG��ycQ�	��Q�s�|�M[Bh��/:J��WN��Pv�ti�����s�~���[�Ț�{����Y�!�AOe�mG�%����U;W ��kGCL�+>�'`�v�Kh9n�x1��U�P�67z�#��}��^nA��>"�޹��>B0�ɜ�Чay���Wj~:��M�ƭ��'�+��f�O��M�?pƎ�u�q#V]/�H$��i��3��;ps�F_A��$c�q@Y��}��ui���Vaf��I^�J�BK%>FE�F������Z5Pux���Hթ#�Ƀ�����m�)_��}4m��0�An���m6#R����B�T���ԟ�uqQ��>[
W\�9 );�90v��w%?�2�?�@�
鶪�%)e�J���8}m���i@������T�����,�`�^.� u�_�5[�'-��>�Ҁ�$>8&G��lP��f���a�j���@��-��76���7yخ���9�&\�$4eR���g����� �$�qS��I�oV���=��t��T-#!6͌DS}�QX�Ls]�V������%��q%ϗ�5��EF��y�wF��C��O}-�ٸ�M!Xę(YwbL����ܬ"W��F�~�NAh�HI?�; �gE���5��d��(�n�d��h�;��N��_A�A��m�[�R̘yk`�wm�����Oɭ�x��he�c��A���o[_��}�l�v���>=��l({����gc�;��K0�u��B��O��f����9�*�
x��(�@�N�ã��YJ`���p7��}�ə�� ŵ��Fv���V�wbq ?�p��6�B���6�wPy]�t�Ζ3�nc`���\��EB�����	��2��P@zx���Nx���3%2���A)s��'^|�7#pH��1W|�����l�0��A��?�=4�Č�Bd.��)�/:�	,H,EQ���jvnh*'
�;;���	9I�V�kdg�|#bbׇQ�[ox v��0Y��8��3��N;�o��aH,��߸�>ڐ���B��wv�[Vz,Ő�8�hK{�8�cM���-K���"�����T@@�;����(��D��ɥ����v�@�胭�B� ���`B���/K����Օ\
>{Y����c����C�R����-Oc��q~��M_q��c=�]藷@�t=@y��b!���\R>���"�i�Α��3ݧ6Z��CZÓ8F0@T2H�L�M���f����W�|�翨�)ɪm6d�����lpw��dc�v�v��8V4 �/]?�3)�����U9��H���������z��l*�ѓq o#yؒ�3��wlX�a$nKt��j�v�Ʈ_�:��!,o�q��N�}�mʴ�f���O�f�^<����&�Ԫ�w�"�L�];�%"���|�x�?O%�H�fumK �����d�ќ~B�eytJ�� �XQ���)��N?���	�c蕷���g�U����᪞x�F�Ě����'�vӤ3q��x��%�{�"�vU���Mz5�ͷmy�s��' #��`��_X,�F���>홡���<9�H�X��V/^�qZ䒖6��^S�e��پ��~�x��g���'�ͻ�����վ 3K6E�Xa�@���lj�Zu{��������G��^�軪�Qt�^���+0��iGK&��;G2�>q�����r���Bd�,��1И�;M���ͭI�f.��U�e���V	n>7˄�������{��m�!���d�.,���6��^O�M���1�������]�[��7�w��:��ߏ��kX�fT��0({UQ�����90/�N]�/�@&����r�_:J����g��!�'O`\Ρp	������&�{u:u2�;q� �}�4���\&��!_L��h��A��^\9��Iʢ��P3��;T�=(���S��2r�$��q���J覇��춱9DL�Q��A���J�$������l�$yP	�>�yn_U9���E`�������p+[w����/u:�/roY�rj��G�@��t����:l��M�-3H���x-d.�?:E���F�
�V92��n��U����_cH
їK�og�uf���ZAe!�X*���f ꉁcw�6�M���ˣL�O�Y�z�	G��eP�
{�S5�2�CfZ����FRłG���1�j]��}'(��93V�)�/{n}F��
~\q̏��\F�l�;Sl���z�g������:�9s�v)���Q�Mͣ��>��\�����|6](/�ƿ����ę[�2�90kӤ������{���TJ��Y��,_,l�e,����;
��@ܤe�z�@]���/k��_ ��\>X&DߖWmZx���Z�%�w-�#�����n\.�b�-�pڨ���C�W��q�Ǿ�s bg��/{<��n7*�7n�9�-"�Rn���s��s���i�������q[�!�)����9ö3�\C ����|��n��y.�����]�����m`y��N1&(EX�ar��u�
JpRP�x}G��8���fE޼��AfD��i(z�\F���7х�z�4J��
ҙC�X�,WU�Z�\��'�k����[�ұXGͮ���3QI�P3F�E�O�"�V���:�<ޮ��
�Զ6L�f\Z�ݷa��Jw]�U�S��[V�&w��쉖��73��>�)+���UR˙0�����6�VCIôN�)˘���]�jK��Ae�}+�~���~-��@�,��[��������F�� j_7��wU�hQ��2;��h��T �"m�r=H!�MY��~{��Dw�����qH����<�X�V��3��Sh	�A�,[(QIPZ�}��_�Q����fv]��p����;�>O��l�r���� i6���*ɸI��x0K���'�#vL*,������ �����k���oi!�[gVA�0��q���[Z�TJU�y�3w]��;�,��^�8�e�k|�Z6���ɶm�H�Xz��=�%p��BF�h�
������r���E���_ B�"�0��T��5����C�m길��􇡙��(pD�x�b+cX�E�祍�rVĿ��l���.�Z��
��?��fw�ǘ�:P��2�h4�� ��9�{�!��� (�:�4BY���sH�B�z���f_���ރ�w.b�@}%���S�o�n��v)��:� Ǉ*����B3I0tx��l�oO���v�Z��.�D��z�</~��A��wk����,Ζ�iG��WgЉ��R��MY(j w���]��o�"%�L���%��}Dl��	��=_ɦ��"��̧D�o�yQ�[�~ɼ�`O ���3�M��Z��t^�����u��k�J�WJo����A�e�K\+����[������s��[ .�3�t��L1�~!o�j�'��f�?1*��dd}�S��A�����A�%��Gj���x��M1̘�QoA�Ա��ڕs����&}|l�ϋ�0�,��>��"�z�kP���q��K"�1}l8Ld��D�o���7�E{��dS��uAC���T��LV8W4��V�����i��y*,��e�H�]@p9!uE���"��gfP��Tu����@&�!L��q/�~F���\`�Е�(��]�?ۣ�����`0*.���O/b勇 4����[偍�FL[�r:Y�Q�����@�c��h���W�"o��>P�c 'nގO�NL�Av���hE�Y�r�b���'+���n�A0��HN�C(�B;��t/���L����_*B�Fe�½ƲaA�>HсU�hsJa�<&�����G���$Xi��F������scP�w[2w�����4䨶�w��.zf���
�����7��X�(lm����{�3������۾�7���$9*���.�dA�٬�9��໗��E�e�����*( ��[��߼w��y{�����L1�����k_5C�� A�?:럼p@S����*3�A�٘q�p��<z��s�q+���[��%����h@9��R0����3�!��8���+}��z::��FV�B��6�q��&\�T7_��ʷ�]���^N�%�x�����~�EkJ��|��`	�����������2��7�s�3��b�J6��)ש��P�����KО�S+�g՘�I��
�� �:�9mAo�ʹ<�����@���$a�\<W-�]���?b�9�(���:�O�K���e���v�|���EDc��1:�j^����G�OJ!��`莉ƨ������>����t>t�W�V���mb�&�W�y��h��Z+1���ZO��bW�h�C��;�MF&�Pdy�b�*=,���1���)�'a8��	?�]�)�p���?t�@ϻ�d;���Q���@�s ofb[e��QdÌ�r�s*�ie��}6eZ7Z�\��{�Ś}W�+ :�[��dH
K$�����e.����߽0_`=x��;���˗

�m�'ܦs�_���.���k��ю?ǅ7�
�ǚ�׏�V��	�ĐMc�6������؇b�P^] |�@��:���dA�I�T�-F�%\�����0x��n�}1M�����*���QpNP㩍����i�%�f�P�U���˴�$p��2��\�KT9��'�������%It��<9+E�����`�en�]�K[C���T&ؽ�,АhF|��-b׍�d#���!]A#��7H�L��&I[�*�D�h_��!������ՒoT��FV����A >�ƺy��ڇ��EXY�6L�*y����o3�v�[��ZL ـ}p��l_��J� 1c���*s�-%UK��U=���[
�����X�i*�%�|���)X�|PŽx��
!�}=�l8��zN�Ο��R���W+��+��-ljA��pQElҩ@=��V�����jMUo�F<�.���^H++�%�( �S (vT��7�؆���&c�ߤ㊢�s��,ֻ=�S��h���?oxC��"8�����g�nϪ]Q�dR���2m�6"��w��Z
�:��*�X��wlן�7�(BV$�=��)�nX=}Ra9h�&��u]Wp3M���I�ap�l#���b�1Ayg�����/С�*(��/WC~��9�ן��q�.U:��s��"���v��>�>�����qݔB�M�}F{k�7*�"��˶27�Z��Sl��ʣb�qXK즮��e*Ya����#&g�g�%�zo�d�8�>�T�>z�����;w.׸)�LB�n�j����2�u6ݯ�FO��7z~��
�����	��
:f�W6��)�J�yC�U/���Ƕ�-�b���v�����3o�T���h=FQ]K:���7��7T~'�3���φ�Rd��˚D��,�G�����b�Xqy��C��3h �9g�\ED�ə��%����J��j�jڲ�Q��^��=%��	�%�B�s���y��Jx� ���nU���z��dE$a�/�
Z�:�� V�Na��ª�[����?o(KH�`���L����+l5U�┇3j&2����o��i����nBT�qZH�{�M S��R��?j����s\�	U��_�}Ӏ@�۴�E>�uc�B
I�u�$&�<O��KD�U���_���+� �H#ߎ1�mL�S�^:+���;��V��]͑�m��A�9��jҹ?�i%�Nb2Lof'��ǀ}�Q&�o~����E�!�RZ2�%�i٘7��g[]��Svf	�J�7�}d��0�>�m}KJ��̾
�솻�1j�Pfy��p�~*=;�0�Κ�C�Zf}���36��j���:��(�>��n�T�U ��fS�j$�U4IZn�`��y��+�N���L�%@�g�K�OY)�a��uc10ā�m��ߵ��5�t��&c4��XQ�3������p_��NBs��n�s,X^��+A������e�������o����ґg�J�� ��AO!2�g�L�+�\�ZEl�����!�[��Zn�So�G1娂V{��|�%���Q��D�
��Fm0��z_�y9�+�$a��T���7���YCܔ�fr�����H��?RW&7�d�O�J�"	{���!v�/K��s-�m�K������SxhgH��Q�'L��l�ҍ9P�E&��#�@���y���1�St�(J�DO�����G�4?�� 1ї�s$k�ѽʟ{�D3aiAW��s�Y�ˉ2׻k@�n��L���=�������Y0f�pQ�HVIҧ�iT�u�uA���z��#���|�Cy�_o6k��]��v��v�� βc�,��ԋ}#�Z:Rp�2- _�`ϊk�u,�K��w�u���3��~�b&Ci�������޻&��J�>:�p����J�5�+�!8�0�2?B��h�#jg3�2�Ў\�r)+�jx#g �q8'��F���JkV�+%gZ�Ӫ`m8M���x�`�/$-Ѵ���1�~P��n--�d?�ݿQ���X?��M\��V�?���� �:D�Bmzi������<�ԁ_�%7�r�x���j�@-U���}��CG��A�{Uz� y(g@��1�2��]W��[�J�9Yz�
��e�`:~����f��j܋a�z�()c�@��EA���[;_9��Z����Q�5A`�uk��n%�sV�Uυ�B1�RcW	)%H�w��a���T�4Q���O^V �T��N�_���� 5?���Z#�
J���wZe�!?
S���1�������L���'~{h��/�^�W����1;��y�mV�=3�0a[�H��N�IbS�k0�,t���f���ڮ
8F��ڟ��X����F�1��B�,6|�#��'�5���"��S�_�x�6:���Q-}��jx&��M�hK"F�܈������:����]�c&W��O"t�^y��jG$RKr��|q�����������,���VC<[�IU�دī۠��mֵ� ���`��Ј��O� �8��z��mDrn��yؑ� �r<�i�k�Y�i`:�$O@5~�f�*F�w�bJI�LC�C�/om�l"�j'�!��v˯�he��\�.���<My�����b�]��=Rŝ	��礂���2Gy��A렳cTL	p(���K�z������J��-�n�'X���oV����VpP�����AK�	���B�>���;<�-Kz�3&��ڴ����͇ -x�Ȅ�yYe ��j4Fs��w���Lz6��i�\��� �Gu���Q
�՞�������v��#�vƁS�OD��s���]*`Wp;�a��c�7DA;tו<
iٖ@l�,S�2�=��Ū�-�݋A�h��Fמmt]�>�ıp{d�g	��4*� =�D�M,׫s �މO ��
�»������,�.�H�O�I�bg����S>Y�����_d��.9���B �*��&%?�F:�w�!D8���j"��ZK�n���
+���ɺ�u[�2�nq�Z��0҃8�qS�cQ� �M;J�*��Z��i}�sl(�Nխ.纒��9l�ѿ��� ���v��m�?i���J/�W�����TV�����gQ9�hlJ���mhm�f~�)?�'U�N��6I�CT���e��ئ��ճ�D�
[� ,��y�(�e|N��j��ƨn����h�>C@Ô���'�|�z��-����4���%��´T�;q);ҟ�������n��3�Y%��`�2хLЧ��w��R[
��s���yW�-v�{�u�����S�D��Je�D=K�y��8�S�왔集����Xz1�WJ�de�/B�j1e��^9��e[��|�\#]���3�v1�wBQ�-��E-;%�x5H�7\�ΐuW�O8�*V�kې�̶���4�<d�@
��}?����[�1���<q,.e���2<�J�1}����S��G�ܯ ����lV����\�4��[8��+tq�M���M���Y$Qؐ
ߝUV6s�*���h	M���ۜ��B���6������^���=^� ��6m�Zr�i�A�;�ӕ�,�Q����r�ɠ�OZ��B1���_n5�F&ծ3J�tb��i�8 �E(nÅ�J��;�h=�ȆS���P� �=��u���6b��>BRK��WtK۱�)d�`ڕh_���"�%�.�no���D�FJn�r�<$��'���^���6�Qb:�k�a��G���W������2(Ϲ�10r�VX+��NVۙw��d�Òq��a0�fW�,o+%-I�/~<G�B��u{�f�m��h�ڞ�}Qʛ9�7��[]�&;{h�Y"��d���yfS��6X�$6�F=K����gvT ������ ݘ|f����࢑��b r��[z���{���ҍ��0>�xaD�+���}i	�q� ��nQ��C�C����a�ފ @��3~�􎭊��Sm����}y�ݮ�^�I�������=S�	�P�t T
=YV��{�f�t��e�F��R٠�5���c�9I�Ŷ?�����H�Ju5c�0BVúG`-��d7�ͅx�c|}f��U� xHJc �-�<�2����(<B,*ς824��G�"�1��9����59څ����8��_$=r���ԵV�8�W����ʠL]s�'�b��:��qfW#d�w��d]C{#�I=�@��G8<��� ����43'�����1z�Pd�$�"=���q~�Ҵ���|�YQj���rw��&M�ܶ�N���I�ݧ��Xr�˞,BQ��	[|ď��d��
m�vR/1�TV�fj�K��^07�;�/�<΋K����U���`���Ç��>�����@|�Wi�x�4�Q��f�LmByp�ܫ�����y��Ⱥ1���֦����Si��NY�A6p�Z�M�����J;���u�1zN��l�9��N���e��$�+�? ��/�����a��򏲲�`�R��v��:y˴8l��p;���L^�ª��2{<a��G-������!�*<2M�����^{�+������6����P��ʩ7ƹ���O�Rs�̋�� _g�"���~+�y��wL������9���%��G���lC�%���ӻk�)��)��ڻbF��G��{�8���l�{K��ç�K����<�DK	�|�ٌ���Ay�[�x*�Ir��Z��UeC%����|'iI
o/yX d��	�}
�����,!y���_"ޅeS�ɦ����{��&R�>8�T;� �!q�X��&��Њ|�ˌ�zʽ|d�Ar����.Ұ�B����u����� �hH�����o��+���m�X���5�0.&0�D���S8Zr��v�"M ��T$:��~�tE<h����
���)toy�����j_�p�Nj�dav5��eq4��@���6��y{�7�	�,���C����ӕ�Y���alC�sg��H8�M6WWؼ����bG�bm���$T���x!sbymC��� #��+������ T���:��j���MO�%�-X�^�x����a-�c��D\.9�ѫ���Z�E�ۚ_{��B�%W��P�1�A���6�����Ipa��eX���ٷ�T|d���7]k&�05.t���crUu��r�,�a
�V�!�`�^MG���F��fF\݃�^]-e�)�2j=[Z�t=L�+,Gr�a�&�Ϣv��m���s��"�37�bhG�ؙ��9#����0�"�^O��������\2����^�B|��LA�^"�U��wh"
����t�����2?��U�����-7��0��� �����b��=S�Ɂ�*@`��}��!%Zj2x�xd��T"$�H� ]+A��n���a���
�_��W���� 7;&V�*�D�����G��r$�X�h'�j��lb�H8B/�x������٘$�͕�>e#
P�����W�����R�����UT���[�E��b��&�f�q#���;��EE ������r���{����XD�<6>]���AaMC"����FP���Բ���~�Bk�&�݁�1C��SO�b�����y鷔�w�A�Hc����r� \���Q��<ރr6�R2[��c�[#�z�t�?�sIi�_�(�P	Ug@z_�,}���Y}\��7g���2>B���k�g��4K-�]ŌI5OG�k,G�M"���-m��&�3�HO�0�����j$���Ml�"9����V&�P���>6��A���&��w��%@��B�g[�y9?��7�Ɛ�T��	�7��:��+<Zϋ���`�L�~#�����G�j�8���t�T%t�0G�c�&,��}ċ���hp�"�p�f�|а����vRң}!�^���� �Q�QV�������]�}h�1�\mv��'F$H�).^J ���g�X0¤k�T��eqt�:t�7�^�^�����τ~{�H:��\�����=���פV���Y�c���צ2�+��=�r͸�ch���Xu��$��yݿ4c��	g�ß�1a��GWC��͘�zLW�x4Sn���C$ڴ��jE���A������&ZԽLE��^"�~3�K��T����v)�`��l�-]!�Pu�G��n��Ӿ��!��wU�}f�C��v3}�e4��.�_z�����Q�j�JL,��-L�Ɂ`B�{6ҹ��Q���U�A�#��YP[Yh =�r`Db#�̻��K����g�S��J���H�����*>||iy?��� ��M}b�O�cz�I̲����)�]jQ�ؒ�p-�b��h5�i�����\
8Wou�]"z���M�
���t���]�f�F͠�����yPH���$�7�meeEQQ�{� ��%a/s����h��d�
ʫ�u����y!��o�b������l��?���C� ^#�cr���7�0�"5��%?nUw���*KScF���n���P5e�S����*�*sA��qң�6����`�X����S��,/��!N����s��N��%w�����^�)�<����Z�榶�'!H���Ѻ�� +�� �:h�ģ��z(�yG�uX�3�����Z�A>髰�R��,��n�k?�6�"�^p��~��_z�ik��z�ܘ-sa��_w�.DB�G�G�6 �inS���k�ڎd�K�x����͗O�4n���q�i�)"d`����Rq��.I����n8�S��1D���ƞ����.�D��KpM�4.���*0jqT����S�1NUX	h԰����C��C��Ϛ}�� VQ��BN���?�X:l�v�. �Cz�#D}d?�����y�sq�D�ӗu�0#�x����(���T�E[�ԩ�3$����S�G�=4��SsڬV@��ή�{�u�%i�Γt��V�zR"�o�>g����]$��x7��t�8;.�cT����Sq`}�V�eW��ۮ��A+G�n�&����h+��9�&�~_���C`}�[(:�d?��� 0��@�[ޢ��'r��^]?=�6�VN�tۆNKH4=�n߰)' c:#��h�C��B�f7#��Z���59���)o��Df�u_`Q�u)������P�`zI��a��/����5e�n]�X��zZG�6�,�+%h���劙�^�%3z;��W0.��}FcH�p  ��~��Z�7�'ݗ�k5��vJ�&8(,���s�� ��N��_=�RW[	���75���U'�Hq�7q���v�÷��Q����?�g�f����!��Q�AQ�"�Mސb-ع�YY:!\��K͹���
�F/F_">�x���@�}l	=���\�L$h�KρlY�����Y�TO�mM�LA��U�_2E!!q�8�����E�\���Ȉ�A�vیW�9pd6�M�� �	
CV�u6tw�(��% �6�]f���4�{R$=�y�a��wu=���� ������Qf�s65���
�K������t�[i��5�<h�7���G��SA@Z�$�t_m�m�{��pl���E��V��g8V9���܊k��P�}���{�Q~'�ǻ��<9
xJ8~~����l����9���fGNǩ͛�x7B%K
���'�3W��#Ö���*�!�Y�A�t�tOI��D0�Tv
�o͉��ro �?��7�ͷG��ʁ'$B\��|�U�L�1���u�b^��@~&~Z]q�o>�*JhUx��(���ӳ;\sk���)�ɯ�"�{�i�����4�6�/�-i��Q	x���}�=�r��gm9�Y�r��f���̕Ǥ/
^�e���X������#.F�`7mq�M'�L���ȼ,7�i���!���1���-�u�� J�^1�1��"ԉ���͞�
���>m��|�3� m�s�M����<«Vy���B��_�1\�6xh�&nQȱ4�����.p]�����N���@!�=&lRYHݥ[,�V܂�/P�OB/6��;��	��c؈��EN�?�rA ���؝v����E�Wl�,~z��������.����:�b����N��1M��6���fs��<�y�E��^�Fxu���r����ƺ���m���ax(G�uD�3��G<c�Ar{�6�Ȼi�����'�M�:�����"~^؏-��110�s��f�0�(�Sz|o�XON��.Wi��ע�Yoh�G2�S�ykta���� ʉQ�Q{�,0���j���ʻ��<��i��OwH󥲣��Sէ���������*9/s�LbX���X��9��� ��x��@���m��)��Z]eE�+�y�}U_K���L����+ٷ}�ɔ��-��KO��xxq�S�@�P�tY(��*�[��R4�OE�P`��_��/��H�W{5���}	�T�TD�;��f��k��%b��q^�l���h�^������Mbށ}��IH��i��c�+��@G����~.x*q���J��2&r������3c8%���y�]b��Ŋ���/Z�v&��@����eO��th�O��y��`̛7�uYZ��i�#�K��ʆ�F]"�1��@�\eA�Ě@Z���֯��ʻI�^�:qGQ�ܽ��U�o�{s�U&v'Q�A�T4�}ݔ�S����$w4�Wi�����-;"��G��p� ��#Y�>=	6����ܖ3�o�?�ƕ?5����ݡ׺u9鬃&Z���pcd3�2Ŗ��5ȁ�8:��>�W�F��[�`�4���z
]k4�ՕJ�c��xQi�r6vz$�V������P���c͐�̨#c���?� ]�%�n�(Ǚ���J<KS0lۭ�;"cH���O�Xw����M�M���Y�)6�{��;���Ⱦn���@g�1�j��x��g�lB�,Pmh���6�&8UW.���q��'R�o�spk����� مhY�^�'KX��~)��/�g�"��ٙ���-P�����e��,��&=�>ո��@!��`�L�7�q�����--�%�����
	wL�'Tfc��qc\f�rN�~��M��[���l�H��Q�P07�E�w� �`u�6�~�9�~�oyLH�qe��ŀ����1QyJ"r�k��f���D�aqݪ^bx�͌�Ja�!7ڜ����O��h�D܁K}�����`g�W��>�cN�nō���.���C��W_�J��i��K�VnHP�?�6�겷����k뇈Y��L��T'g�T��6���b�([��م�p{�<��;�-�o��9�Ҷ�;+`>��v�n��_���a�irq�9W���++2��'L%�@y�I�|�p>���aa��C?��P���W��Eȫ�K0{	jg�5��C�(CLֈ� Bs�-` �s�C��f� �jb�.�D/0���S��9ܖh�S�S�w�=U���L�dH�V��4�8�۲Zˏ���¦�u�͍�9Ұ��K1J¢{�=~����[FQ�����ǋR0%1Mu�	�plU����	��l�Hw�O�s�EVf�h���
�'�9��� �+�2\����/t�P�oݕD��x_@c���q��	�DL�H�p�凎�j<�i��ibگe���a��C�~����\�t�bi̒K��X�0eᵗ6��&т�hS*���^mz�E-����/;�,G&D�rZ~��ԃn�"�×v�_?�Fjӟ�WG����jz�v������ر� Or�-ݱ!�1��.�\DOZ/pJy��0/5��N��ǵ��S���yF��>�%d�R�E�Đl��*�D���
,$j	�G��J�#���X��A6�1���x�s��7�4�@G�ux���c�ʔ�x!��Z2t�����!AGk�)�J�\�ps\�p��L��.?�cq�ͳ \�F��R Fa�.���y9`%��d��r���K(s����dB���8B���l�Ǘ!@��ӕ���̛��u�i0��Sp������7��8u|{�C2:�`���a�u��*��xV�d�+'����9k�?"]v��7���1�t�������%S�� ��ٝI��*hKp�N�����D/��S���g6��������9�>�T#���iN+�X&��;�C�仌B�� 		�0,-�q�AR1����YMU���9�c� �R�0��k|�d�}��S�Y����\�9%��`�`xɈU���R&C�I=؍x=0���.{�v���b_���� ;�emG���2�L@�F�p�&#�8K�
)v��dU&�	m���{u��W�ⓋkL��:�|#�ZM'�S��z�g�\-!��I�W50���u��al�}�w�sX�)�1�[x�Ƞ!�=@�[<E�@{1�b�zl}�s	Z|��c�B�H�S;�`���K�h4�w/Ԁ��H���������I$J�s�m�:ʛ�oY0�)�)-�H�`��݄�	���:0U�骹�y�Wr�5��%�0���@۵ ����9v���<�n�,�}�[�p�C��jD�����d��;���
��~V�R�ٷ9nL���C���B}�������A8eK�~��3�nN�H����,�s�exG=����ޛx��|�n`����*H����-$�	pa>8����=ଧ��8�_ ��T+�3%�������z����)ɴJY�P��Q7;b1�A��,Α�>�5�P�ɖ��]��Bh7�=�ZKh��&O$>|�pSH�C��Zȫ� 	=�6M��GH��{�M���۞S2��=���A��a�������S<ּ��e���=�p�}�9��lO�r7z�Yp��ʂ��+�^z�[�kdlѯFB赏�����G*J����<n��sd#�S���H����5�+������aM�E`*o�lsͤ6�=0�����o*�-R,e�9/� ��qM���{)�{U��e�s��d���̸���6�[EA�r	G�wN_
���V��TF7�Z�@�]���'d�x�>���
�o|���W��������PAdT�a���i^�W 2�qV���'���1�Ț>�NCiU�Y��~��;�����A"��F^�.&�I����]=@�g;/ �+R;J��Ra�j�W��ۘ4�vY{�� �Ͽ.�]$������##P���y�:z��B����.;�.�2�{���AV�Vmj��_�(`,3fc^5 ��Q~��{���J��T��o6�\]!{f$Lض_P����Fr�SA��)�aĭS%�q����@Aă�t�S�k������!�PX���	ʃ&�y�;�K���-�X�n
~��mZp�Ε�I���nwC�+���� �p����D�3�{��N���NԈc�d�	Ԫ�y���坾Z�74�Лl��U� ��E@�N^���"�$�{6�r���Z�Y啖�@����\�Us���F�ۅ],��^�������(M�A���73Y^�`7������(Kj8C]w�b����Z8wJb��B��})w�[B���U\2�P^~4�VTֵ��{�%��r%p��:��'U͹��,�U�L|t�0�S	�5'pޚ��- �%wv,�	�_������\��z�N����ZszH薓 wv�^��h%��S��%/13�V����J<K���v��u5"H،����"w��lz-�`i���=Sf2S���Z|��a�2}�%x����.ȇSG@���5#+�h�Yvc��m�ͱn R4A�3#hjκ��6�gܣ�}Z����*R��1���T3��7w<��4�^�3�3��X�����h��h>.g�	�Pw�/��數���/*`�.����1b���g��oF��z�"�ˏ��N���:�?�"�����6>A�O�`��fJ��Q�b��c8r�:��>�i�I�� �k�Xo���d���`�j-�%k�U�޵ pB��AB���	��(���;�.�3L�y3�����vy�FuW4��iP�=��%K瓎 ��c4o�����]:l�]4��^��<�uZˉ3�~�(La�4�e6H���5����s8\�jd��M�z���KLX�b����1l�[�7�:Y~�;���˳Z�'����ht�_�_�x�hM�@B�E-܁Σ.�^IA�*�m�e�G������Vo�0o�X����v�Bu�jE�=7�ekY�1u�*
����.��X�O���P�&=���R`;�&�5� �T6�����H�&ri�@�n[F/��8� )p-�Q���x���]�������!%���$��4����b�Y�7vH�?��?������?E����:�Y�K҈uD�����͎�i>�aZ��/�_���\�������y�l]ֿ��-yߘ�H�VD�������H3.I 
�g�h3� ���C�dH�l�mQd�@������}~��ri�G�0�x�I��4�'%)M�XW�@fO�.co�q̇��ԙ���@d�8�.�K���j� tDP3sؕ~i0�m<���!���ϯ.���i�}W;�x.��qs.7�Jɀ�U�K�Kɔ~ː���߂6$|~"g�D�tQx'�e}y�y�/���8$㯚}t�E�,�[���w��6���gK���v��\)�7������2����)N5$>� X����*�	��n/�T��=Ԣ�-�NA�u~�90c�jꄭ^j*��.�$?�[U`O"���_G�n����n4�o:�؅$Xk�n,��6�0���#ƙ/�+���]k|��T��!Z��`�B**z�҅�)���������[�<���P&�t@))s�Dr�1b�+N±_�E�Ym���އ�&�����J��oČ�U-���Ϛ9�t�����Ο�j���}��|�����yh��7sk����VC���v(V�X�D�	�������qS��`�_��̬�Uo�m�lJV���F1�T�t����\�ڛ���sF9�������nە�S�d�r՜EޭTB�|�!�*p�C���3C$���k���a�:�,�@����(�O�1���ࠔ��/�QF)��6���q�W1TCj�O�F��!I���1+:?&���LtV��&�#�V~B��H����>�.�
�̗�)DB]�)��#�qJ�P]$��(l����j����VЃ�R�y1��@j�Q��������
�5�<��G]�tؿ̏��P\�>쒘g)�K�P�X�`Q�Z���U��tXn�Tbq���� ��ل��Tc~��m���Q�B�+�+�4k������)����Q:�unϭ�2�� JTYZM5Z�B�D&���ou�nd���P��,��;��7�L�������c��C U�R�Nx)��Т��g��
m����Q�SLX���%�%�[~ǈ�o�	tW��ʰm�o�C�~s��#�A��u�
��F^e���v�yE����K����!�y���WO�z�U�m�oX�8�]�<<D9�:����>D���!1���V��'y!�Bg���̗��f
տ�*;i(M��U`_{y��K�*��UXzg3�����-�����ME�`��P^��0�@�
�h���E���<�s�xkɨU���Uͼ��SʴLc�P�i�,5e�E�n���%gw!��z*��M�`g�.'�A��a��
Q��g�H���徛�ss�c�7�`��ް�AV�Y�l?�[L���b�� ;y�*�H"ľ�K�<��3=�������$�-��n9W$o2�	ŞO�0�T��9]��$.*̓��J7�;L�(��w����@�l�wN�$����!x�#�@�x�ې�i�3��h!�P8�sH�}��,yU����S!􊂫�hD�^��r�$�4?i<n8)֥�_��E"�N��.���)d�M��n�H�����eCL��u�x4�Y��
����Ǚ�ޠ�t�~�P��UR�S��I�)�h֫��R�v;c�J1P���:�e�ZS}�j5��<[�
������\�+(��}��J��lo/,�]�8�^8%Q����F�jM1�q�Q��M�	ׁY�g�:27�Nh��E��{-Fۤ��~e_|Z��sӐUp�,c¯��swϐ�b^^�tq�H���֎g��;e��Dt�j�ba��^�Ҝyđ㨛�Z�j�N���ke�w{��qPac�W�Y��q`Z��wK��ղ����*S��X�+և*x�߾rEj~�P�&�.o�&�ʾ�w�^�O ɥ{D�r�ẵmuj���V���pTp/��7��\}}��7�i�%�c٪�l������4����Oڏ.2�m����W��B��[��5(�~[�[�`J�r�������J�b�ӧF�)o6o���$���N5�=?�C;Y�.�dX������˦��uI�R�R��FI>;{�Y�S�L`���V湜M��0�����S&n�D)I仰�ι{��[� M��{�k�EK!��?��-l3i��:&]2+�C8�<�C�7L���0&�̃�R��2Y�_��KB$S��u}����`���AB�Bk��N.vB������� Q��������Ȭm��Bu�,��4Ae�����G�-`���g��R�(9枺��	��R �0�1�~ƚ��b%�T'�s�RgT�{��z�a�v�P�Pg��%7y~����g���O�"0����F�����.�iT~��av����bJ�L���Ȱim��OŶEj����6�B��<t\�I��J3e[d@<z��1��?�E<��k��6�{�Ϝ��L�E\\m5����z6֐:�[=yh���@���;���v�~%��URT�KD9��qn�62�=EGP�#��X�5�(2!$���fR�l�&B�q���a�dޙ�<�ۆ�"�>�̓j��͵��+��G#��I�n���8�x�˕f�F��C��ա�I�bj��Q���A>�W]�@�ҩ,��z[�Yd��P�Ǵ��n&����9v��T�ɲw>[��.�p�|��aH9is_�d���e��@�t�I4Ia��/#������5�>q�zz%����M�P�z���z)��+q�~	��^��)\����Q64�K�f�Y(��?�W���!��/����ƠE�J~y=4�#?Y��:`x�<�~r'��d5�w\�щ�a�
�5����"�2�~�PE�g�!�Ѵb��|J���/�׽Q�O9y`Y�C��ǹ��7��_z��"zrc�y4./j"�$�π"l��<��\hqS�	�	�*g5y��J��%Y#Y�����y�����.E+I�&��N�ݭ\X`0v����������DBVK�>�J��?08��1C���m������^��m(�nkGȃ��&O��2dȲȝU�GĪv\eUX��AZṅ�k�(��:�h�<����l	�aF��+��~�/e��������Ｅ�����ʙ���-�����Iq>����+�$�3���sPwb�џ��6�����͉�W8�1\�p����M��j��9_�5*�?��)�1T�[B%����Ě?[\IБݭ��g���}�m���~�Pk+��k0��#R���e݉�7���gnL�������� R��RQ��gλ���ϵ�g��8��c�*�,zr���f���`P�f�	�ך$�;ʰ��8��C*t�F[��0ȆGFmC�nVݕ����&%lr$�a�Ê�-���⎫Ӣ�O"]���Ue��z�C�BCv���������Ly/�4��h�0��/ɠs�'kR��ᡈ��f�{bc�kK��  ����ɘ���O�fُ<�$/��@˽�_�~�����o��ڸE#���\&#ݿF7ew�G��H�D#'�H3ؓc�;��`q��k�����Y�e5?�9m�JP�|��e]��+��"���,���l����
���K~z�U�̍�t�6w��r�	ڝ@��D�|#E�('�aIl�Ίk�}�U��ȋ,�꡺����6�B<�90T]?�
M�{.�����Djr�=�޴�ޥ ��Nf����Q���%��h�:}��q�͌��w���C��{�����w�$�7��2�)O^��Gs4�m�mZ����\���X��S����u0��y�X��[�~�G6�d���p��)on��&�hk��O5���t�Ħ��>p��톧�7����ˇ�:���:��o�e�~��wh���bm�Q���W9ۈJO�><�oX��-�ӄ��I1g��<.�Qk1�H<����x��Ò�����	�����`�Z�ҙ����{�I�7��LŶR��D�d8F 3���X��yj��Ɇ�<�U�W1��:��|\U2��i�C3L�/La�5@��x��������%��.'M,Al����&�k�1wȩ�F���MD."�pB����1��TV�PѤ���`��v��� \���Ϫ�K��`�jl?��jY���ρ� �ah�Y-+PӖ�M���Ze?�C��+0jZV� 0��_����~6+�3�u3��d�m�������hV���c�~��f3��╓i�G����t��y�W#J,���F��֝>�ٟ�yq���[Ae����"���t�q������8ĉh�h�G]k���d��x��#�P$�a+����C��u��or"bި��u ���}]�8z��)���Rl~�
)麉�wc_h��UR�<�<�'+���	�}�&VT|W?���7��j1$�Lj��
3�֝��Ѿ�.�?��^��#[�`�K��x'�!�|��3S8<�[R����<(*hO1]��F�ˆ�^	�u�m�a?����Yj��z��LP�$$ڒ8;�Bp��O��H%��֐$l����B�α���y`��w�������ks^��j�n�#��ozMS˵�S*�R0M$T�z�ԸJ:��Z�p50a��Ƒ@����i����I�bE �1y�u�obQҌ�v�#qw�X�%,��Aҽ�:
�d����M������p[��ap����z�	j�9�x��(=VeI�R�3��c#�F	���B���32p��IBVK�V��4P;����?Ͱ��w�԰cp	(�P�o����&=�7B�4�Z�@>y��᪲<T���Ga�3H$<pi{O�,Z汥�3�91�k����rD�2���x!�S1ͷ��!U��V�:mk
��6`3��� ��#n�=G�U�Ȱj�/�H��V�k1�Y֛��QhPK��K0����E����3t���͒��8���s^�] �n��j�&����CDy�sU�t7��r�C��=5d�߽- (�Xyv|��_���y���.A����)�=��$��{��F���d���n�Cs�J-Y�Jй��Z��u��f�C)�L�6x�)L�[���K�aYS�%�yQ,�{��3=:�>���s�0�rBm�p�����%���.��X7�ҁ�V����:�ia����<ֹ'q73S����W�8�Ɂ����#O	n-�D �4<�YhM��Y5Ơ4��w?b� #gu~����	�j� �[�t{�<X�qU4���/lCe�%��,��O�;>�F�p���A�'���V]}��3`)�y�m�l�?��΋�%F��E�-r
��a�o_U�6ȷ-E�~]��rp����r���b�g
��	G[l,c'9N3`�(%��4�=��&/���!�(_�Z����U����F�gq�X|�f���#�d��"���(�b��|��� dD�����h�,�s��\Bb�����yF� ��{�]�D��h[�e�@�Zq��SbtiV�z�!4��<v� }���9X���*?"���2�r�ęԗ�q����[����(����*j�^�vc/Й]ƭ�,1� i�~ "`7pW�bz��vCK����3���l����&����C�%mWR��D"q������䙝�y
0�i�q���q��X ��s��W����[�t`Lʦ����Ż'�V�k�QX�*����a�h��g�� L���W)O$h���^��=�<��\[
+��cH���x�Q(f{:���<���ڕ���e�B��I"O`���!�Z�A��Y��!�/ޚK��;����� /mc�_9ϔ�{@be;/��0��R����k�]k��,R��m�(&�*�6��_�q�R.�{�'�*�|5k�K�.J��^k%�a�W�l_\ͪ���G�m�}:���:9S���r�!a��뼱�'�Vq�_�$iM94�E��~���ev��|�|bJl獻U#���tX�9��5�=�_2I�1�9 w��.���^��τ	 �M�������p��d^Њ�R.�|⇻�W�|�����;y��
v_9��)հHߪ:7�g�7r[����y\&���=5�sQJ��G�8X�p�D#�� y2��Oj](�IΜL����*�	-\-� O3��a�m@N,�0���QbR4�7Fg��Q{�B�|9xg�r��Ե/�{r:e�;�0a�����碏��b����V��YS������ce�r��n���T��P�^�>�V���L:�<5:Q:�z���qi:8��bvN5P<ׁVAd��oo7�h���;E�#��T�ߣw)J�����&��H���z�'���,&wcɴꨰ��
��P0/ɚ?���U�ղg�R=%)i��6߄fS�R�ST�>�����.�_���{IY����/q�z��a������f���;������-]��ÿT��
��U�hc��Ք��f�u,y2��
wrec��{1�/�� :����X����_�n"�b�ˇ�}�-�.4i-N�����H�^H4P�g�t����	����7NWm������C��A�� ����1���>�Y�#jpL4�V�20��La��6�	U���X硖���=Qÿ�Z1�����ڑ�1z������wÕC�L���q�Q7P��ܭ<	�yGt� CI檫_����Y�H�܎eU\G�#��L��SeC�g�8�U�}��_PR�� *���C,^��:l�\��������z���Û��:� E�qqA1n�?��A����\W�OE���ןjp-���M�E��O΅���`[\M�o�IO�9Y�4S@ޡ�,��^�IWhem����z�3j��hY~�DG˕pp���qJWy��:�?�}��͋z����*�J���,�>�OF�F�F_~�0ac�����ьc�w�^��RO_u�#�9����?��-���������.^&'�<]2>G(\ǆ�3j�6���yh�IP�5�
�k�<c�H8ra4���+�|Ư�.]�����7�KlI	;C��!Xh��Ppb�ZM�X����{.�ـ/TŚ'��v�+�W<t��ʦ���(d���h>ч*�X�X�{zB��?{��PW;��Z��6���#���<�6)�Jj�*��W����� T �4FC�FI�2�{�)0R��	,Ԣ��Π]ߴ͸6�S�N�����yW�]��dA�j�^E�ݿ�*���'iIlV��(iǔ@x'���֝%D�3�B������8v�Ȕ,h��Ե�=f����l���YK����U��&�<��9�sF"t�}��+�5 ̀�&qt�<��MqP+6OQ�}�_�w�`�E�����v�'�,���W�G�0IQP����|$���X.k[µ|���p���C?�kJ%S>-|>�h;�=^�J��K�%���E�h�E�:z��R�!5' h�;h~EُT�Vx��X�����͢�M a�տG��f_}x�����
�,���5�pBlT�hӪ�����>������m�zk+	Xu7ΈoL�g� ���b�k	ဌ���`�P���ECRX:�G�V튎�gEʾ�%6S��h���
��jn���AD�Pf���q�tVu����%�U�y>����:/��z�<�0�.�	�A�߅\am�U�WH.g�4�
����f/��C�NŸ#�\��W�
��>6���x��*����)5!P�vfQ�s����m�`��[�yd�-:��F�����$jͤ���X��Fb�}B����ب��[�?E�����h�
ۂ��*W��s/
X�t}�M���8 ���O3���+��]��ĠS�Ƨa�����8��x�6QH*�G *ß3Ė�2�p�i�����8�?�2���o�)���Q��J7܏+f���]t�(I2���r�WE1c��j��P'��),�f�BU�خB��ߌ���&�a��ߋ��^|���a�#E�Q������_-�5�sd�$"�pq�Z�-�J
�r�b��:M瀡�1B#�Wy7�5d\��$��qP�h/�	m-)�Hz�Gݴ�_���/�/3d4?ݫ�j�񣉘��MMi��5�C:0��5��ags�e�ˬ���u�F����H&įE���qEgi�u�pc.D�I�M�?��Q#�J����^�E�i�*�䌼\��K��N�� ���������sKW��z�p>��<���g!�^鰿ϤF� 
zP��J�#B����W���B��������[4��׾q��F2D�5����E/�7M-�H^��4i��Ө�*"�ͱ�%H�"��!�G&9y����m�������[���S�����H�]+G��RVko�C��������"�ܪ:����I:��<�aצ�2Z	�L�
���Z��.�8�C�x�b�����ƙ2G�E�-����^B���@BĲk��Ԓqx�����9e��Uw�Z�z���[��Cxw%<R�V/�4�g?�ĩ|�H��`�3ݻ
�{{k�5dRY�E��{���ĈFccD=
ւ$0�ԬP�X��ڥߖ5?��M�> n�>������m&05~��U��;\��'^���8Յ��M/;�"蕣�3:��eK�JX�Ԧ|������R�lLd��WZ����X���'��f�4N�P� �E4���0�:B"OJ	���W�nAp�T���1�]���_᠔���7�����(�� We��0�x�6=�?_��_=���3׃a���D5��VAƻy;70}jU#�$��n�)�g�X<�J*���G,P��~y+ɫ����bç�.�U�y�j�w��K����բm�k�/;��.���l)H���T]���}P�(�����O��� \s�c¼]�0H�o�����h�{��Nz�%Џw��O��2�ң�>ڬ��'Q=��U�A���J�g9��[	����U�:�X�XQ�Q/_Asxݻ$�m-}��	��ooJ:��<}&�͇�&(=�zxox>��;�r��Z����͋�{�ڢ�)�[�k���֏�h[�~�����V�z��e���4�]�P�ҏ?f��<@oJG?�'�D����|��Fc�QY8p/h\↜���b�ذ�� �jv��Z$���g��Pe�D�坷����?�v�-������_�t�;h|��ܛ�){��j�K8��u@�����)�����$ ���Sn.gI�@ͬ�H��_J��,���#+�s�_�t��t֡�K���S�����^�x��4��҈���Af*珪e쟐R�y���7���B�5��#��R�4D�JE�Λ�*aˣ�J�(����r�6J��ח֛"�����-��)�7p���ϳ�\yٴ���z1�>��V�ȯѦP(�~!P�ސ�A��0�a��žȠf�ې�G'�y8K=kh���i�Q{?�;)��Ȑ5������������כ�0��#Z4�9��8ȱ���@8b�y��^"5�X�Q�|����֪h�q;�s��%��r4=���2(W��w�=��@�nֹ����wr�,��W�<�ԾN��t��*�����$�e��ٱ���?Yv�XA_1���>�iz���7����Q[M�U~�����u���j)�k���_�|���le3�B�yp���`��y�z*ǯ&B��щ`_��b�G��C ��ܙ~�9��g��x�ț~���#�Q�V�6+��Р� g׸2� ��p_�T��)��'O�_��a��z�h�8���^���O]�v�%�u[KɳQ�ƣdԒ8bg0�Į��w���o,G�9RE��qb�����v��5�_lP�������B�~3�Q 	��Z���U��	Kk��"^�i�X�I�	 �f��MA=2��.y�ѤƟ+���GO� 
I��C�R����V�J���ML�hP�q��}d �|�t��Ҿ[e��!�or���ɞ(�`�6Z��l��ӣF�SD�8��5�T�6��g�mj�О��2�GR����p˹��&G�PΉo����~"]�R[�)�x[=7Z�����z=��'��KC��GS�Ĕ�f����'Fx.��f��jjW�:�	g�О�R����p�����F�T��B�����/���I\P���u�ހ��Qc$�����}Sšx�^!r�_�5AƗ��Qnz�ȠJ�D��� {��j��ƭ���G*�X��M��8�����g@����d�Eď�V�v'���4�:I�zRԘҽv�IA'M1��ˡe̊�_n�w�T�� �77"X"1���-������ȭ	��:;�6XfM�A'\f����T�:F�`R��5
�z�J��v,����d�X���`ʯo@$�E�K�S&!я�TH�T~��!߮a�:�o��@�;5���qrnl��ܦh%N���D{�YkIs����	�?Dq��ݧ:N�G�Pal��@�16������'�T�=�x-��ojC���}^ak�\Q�Gw��w�1`����Z|���-Ed8f!�u�^�i��F�l%�1yl���d��&�����	�{_��*a+�Ʊ��Q�k%?�|�"([Y��2�iQ��vڼ���d�(�qs��A���?��N=; w�3� ������	�c���I
��uID(R)L�v���+�B�Z�r���/3lͭL��;�,�f����w���8=x��]�x��'�T�q��~��AX��=C7T��&�����) ����?'��<R��L{�)��nUXc��7�,z����DœJQI}%�����D�&u����N�F�!��*ʍ�����2޸.�'�W'��!qў^�6�?�}��^+��>T���P�T���'L��l��v ܦ�z�)��!��x���Kjz�H�@vq>�Y��)��hK�dS�Q�hv���L n�E�]Kj|����W��M��D8���_���v2@���:�ڥۊ��Z1JR����׵:��)%�Ū�C|�l�(���$� �&��O��|��6�l	����uE�(L�}���۝U�ш�$��~�V�q]D�J �	�G����E��5q�r��6 m�oY�DV���l�*�P��>��C��f��}��w�k�s�(��1�ߦ�a���u��j�J�<��W~
22�t�s�-5�!�
w ��o�*�]{3���!��-���,�!`Kd��͇gT��9�wP�ߣ�*�:"IuNU5�$aP� 1�u��}軤��8=����>�E��|}'{uަ�~NP�^��ҫ)R��h,o�b���	�_��uE��fh&����[�_��0�k)�^}H�^{<:9ELsj�����S@�����MR�>!yl�-5cV/!^a�s	�nH�^��s<NĂ�%�q��/���ܾ�\�^>Y���1�Pz�&��@ڎ�@��/8��Г��ωa/.	I7�4�wZ��,wϘժt��V�{��+���YN�&��;7�J�� l>k�j�/_pW��^S�]����G�	�.n��o���i��߲ƻ�j8<��=�c�LT�s�>���A���Ew�"�,�؁��{ؤpu�Aihs�1�-�j�A�x�OHc�an���|H�4��͎�(֥�ҐH��>t��N����f�I�I{Қ
ZB!��6w�αǩ�C�i4$��#��Z���K ڬ�6u˒��w35xk�Dˁ5bǕIiɨ�8T��p�y%�:m�����n��� [
͖`�Nm)�P*7/X����-����ӫcCL�v#�B�zP������\�%P�g�f��4�|qOy_G���ѹ΅qh3�B{:����ٷ
�U��_ј�� ���y�w�^���at�I׮:ǀ�iy����m8�j˹�%���=:0�v���n�V���������g��G CNLFy8�44ʑ�a7��i���Y؜?�ɀIi�Q��O%sX\�,�aF:0�+�P$��ƥ-��X�h͓2!Iw۶P=�е�ԭ�c�'�%�p�Yj���'r۷4�X_�a���E���&1B�����kFL�j\��U��_(6�I:ߥ�K��U�/.�i�vh�d� ��a�;�b���{�.����۔Np�OE�U�XP�\V���7Z��mܖQyڜ��85a���>u!�#��&H����q��2�eu�j3El��ة�@~���S����JR��A��]���Ԝ�������߇�J����Re�aMt�5��)��r��K�1U!�f�l,��i���h=�����Ɉ.v;��i����� V�7N�������A��Z�G�!��,�P�zF���'��O8��e�1+`��r{�tv����׶�B�xC��(��g5-���3�:�!܃Y1�r+���]t�X@3�����+1O��"ö�U�(��H�h�U}�2��������Œ�኉� �b<jn�p�qmX�a�h+s&���S�Ji������r*�$��H��`��k��f�����p�֐���	�Pn��,�c����f=��K�J�G�<8[�M��Q9��
)���{�b������6iF�d,�ui��Z�
<��A�B�F�5�u�,W�t$XH�}JEF�}$�մ��b��\!E
���}Ѐ1I-�P1��o�J�*�/e�=/�ƞ�iB?�u�)P��mT�Ed��V��>��/��	��������$�I�Wupc���T3��?�`:���D�T�P�'u*)Q��/��^��f�<o�YO��$�H4���:.,ޠ�u���ɽ��u6[.�QS�wpנD���������	V<^k�Op�q_t��7�wSJ��	�(�w�x�9Lt=�{�%�`�?2���O���iRp_��@�K���$���*)|s"������,5�5/k��
d_������~��B�!W=��L�b�Vy�s��@<FA|�d�<������/�}�O!��p�iW}�Y��ER�⺏���+wg�Ζ�K�����ǡ�� �"+YI5����e<�˼Z�q7\{��]T�#8�)�[���o�������e�4�@�Hfv�S��+{ϩ���{��_��!�����E顓�x�`���_�#o�W���	��p�'ϲ)�!�����(P�� ���V�{g�M���f�)�{����1����:ٔ�z�L4�6P��ߌ<��5�������g}�}^Ps��mU@�ϮY�������Km	͇~����Ϩ�G�'t�nC~m�t�����XC5�2�@vfb��	|/ʁB�=�ک�Cサ
:�l�ܯPzG��\p�\1vP�y��3I(��	Sų�/���v�i�bC�7? n�d���@��~�.��>����w}Ȫ�\1hxQB�d3���@��OFs��:���/��_3ƪ��G���|�y��٧�O�N���)!_��i?>�T�rw�*�\V	�T�mZj�g�d�@�D]�T�!�"P�]�\��Ȍ/���Lڧ5)�T�,���pg4������DĠ�����bo��p�>h1%7�֟��N��r�,k!����sk7Z��8y9W�y7��8���z��W_~�9g�f���C��vT�V��A.4���Ý�����I�W�8��,Am�|�e�N!�Hǜ����nsƜG��:�����4 o�~�?�!������'ק0��Tǿ��7V/����a�����)؞H#T�⭤Q
@���A��Q[�|V�m��n��*���[g�"�h�� ~-�7�P�G���XV����p{�;w�m��o���Uܖu)*�����O�2���eh����
�f��ɝ�R9f]�wy���9�jd_�	��r�{���6���A��������A������tl�K(�.Փ�/ZzE����5�&��o"��8���ό~����z� �w�\�Ǥ��j=��.�����?�R�Rp�=�LϗI��pa�/�C��;�[��p��/Thn�Kg���.7 �~{�.k���	�~#�Y�u�?��ٚՇTBn�`2�P���'@��s�0��[�k�)�x�8��-��_�̎{C`��B~$�)j�hI-���><����z[��D�窇i=�S�aX��c������/P�;�<|��d����-��0�DdL��G��6k2�ׄeH�Ш�nc�֭�1h�U��H�a۳��ʺ!S2����t�Á�W��+���]��~mRA��X���c��|K/��p�[e�_`_���i�p��j6�S��im��_N�	�IyB�e�ڢ|-	:�٭��m�� �U(ʪUt�w
X���2kZ,8.&�}��Fg%�l��Ǹ�1\��fe���g��m ��g�e1x&N0U���~D��V�����t��Z��F�gN��S]��)`��g<��
�&�rmĹ������y���5z �n۟�d�|}��W華d�O��w�X�X�c�+Z����z�r9gO��D��x�􅣭���U:��������&�I���oIt <v��^8>�y���i^'�.��"��ͭN}�XE��鎉\�@�Ѿ�����e������c�W�8eX7��D3Tt���,�~�.��	'�it=�*e`� (Ǉ�Y��,	�("�^^�X脗4e�Ƣ^��3�I��tS���|�S'�2 �dق��.f%�h֍Y�����ʃ��Ქ�aC��ի$��,�_4�,�0�6l�����ޗDs�?�$u����
�����HS 3ޗ�Y5�������0!?B��������8H���@�-ز�o�����qf�sb�͑@��pS���T,��[����(��8\�w{rtRwhƅ�i�����Z��Fyx�O.E��04k��K�!����}�ȭ���KT����snE�����%~ZdT30,)���B�9hC
?,�{ᄖ��(]v��Y���xx|y}�d��>8��鮖��#H�pY<x	D�A�	������@&�=H��qZx5��Мx�
��=܇`� I��9���%a	r)�����Q)���������5٤��,=û\�����fKK��b��J"!��C�Ŷ����l�Q���b��k'BJ�/�f���-�T��L��C��rtR(�!� ���� �smj+,� 526v����R:	:��M��je|�@g*hQ������"�^搖��:�����lF����h�W�"e���P�D��r�N*�����Ά�o����һ�6�p����->�=�Zb��n�tyE��Mj[�L���D�=Ȓ�p�]чފ��>zt�4Pd�ik;a���\�C��}"�ه�r����N�ק>h˽^4�m6���X/c��:��-"�lPa�1�g�dWU���
�#���~q�е�,b,�0�.�q��h���!}��ܛ�S������^������nC�M� ts�/��	c0���n���B�zZ���N�,����m�AP�x+D|b�@�2n`"��o����g�Ki�?���7U�ܷ[�x㕏f�"[`��*W�^3|Ē&����!�p�`����%��M
t�E��W�"��`����j��&E�dsH$��U�o�w7�4�����ќ}��WN��,��?�|�>�=�u[U���V)�O� �
RiB��U���@��I5eCުyĉ�c㧶Z�{�v�-%�Hl'smW��t�އ���IT0����5&�������SJ�j�U��n�^��Q�HV�� i5�c\Dd7ӳ7���QjJ[����9��7P��P��nW	�� Ö��2WW!�X�8A���9r`f�� ��D|��`ZY?Nâ���(���o�;�z���V�X��Q�i�O�V�`;&��0qa�]WCC�����dƒ��|��
�����jk9��"6^�,�Ч)T;g��TLqB���^�%E�����p���L�U��:,��3����H-f?Vɂp�>�3��H��7=n��\�@����ze����̈\k�9L�Z�x�D?�����gc�����w~�Ш��w�/@�NW�TmA��ML����2�r���tD@�^\C�B��OMJ�~�./��FH��ޏn
g1<�������������='�LX��M[�𡗦������̆��T�5RU<2-� �2�@~�$���9F�6~M�W)q/�<�Q���ː�&�|="R�h "�u�HV��DDݧ���1�,���t���H����$׾}w����n���A΍�L�iQ���ጭx���s �h���`9��wQ����<
v�B/޴�Z��Z�(@��űuZ(m8�z���^��ﰿm�O�*������ ��\oD�"��l�k8�O�a]�H]�܁��"���n�w�Ǧ�Mv�����"5�^�d�6(?�3j]���.#I�iVEA�!Q�{`sć}:��
!&���mӰ�Yx�7qWl�R��2N�W+�@(�S$�5� 	���x�����������u��i���Mi���'5B���ӼWQTNt�fc/,,�4�>��_�9�@�������̓��b�9��zk�`�~��2���U�'�x�� JAظtto��UB��Ī*]��@V_/_U���a�l,�҅4�$y���&�lE����!e��� �U�Dz��/�nl�|YCΪ��<��MS-�	Q1j5�0$����b��D���{����h���<�Kn�M�7���N,8� w�s0�	F��0|�.:c��ñGbC�f%���(HΗ��n4�lP��Ә�=����J�lb� ��5s/���.��3漄�p7ݣl*%��t�e
eLac}�x߭�?3� Á��9���鳹GzQ+m�� ����9�<���:�ATq�(n��ɜ�"�{��X��c\��!�|��lisk�E�ќ�t����-�e%�T¹�2`�N�]��Y�Gտ̵�t[��^����3AQ�� �$�"���#�~~�H�d}/y��`?:�&
g��;�"���9
��Do�V��;��Oj�Z1A��!xK��+���*��LS��u 1��C-����67:�M�
}��d[D�W��Q��+�f�umA����'�GU4�RRu[��H_P�F��	��1@`�T ��,Z:(��e�v	b�Iw\���|%�'��cmM9&��\W<ho����\)_DM��@R��6�s�C�V�7!CF�qߖln$��]+���6Û	� �ڌ�$Q�6M�<E�?��,ha�=���	����7cث���G{c�^.�_��$���=@���;��!Y�=9�WH�l�f�@�������:�ȅ�j<�Tk0rb�b�Aj̨, ��W$.mi��z�g����=RQ����G��F��h��!?�ʐ��v)S:�c��d��`ۍE�P��vv|��F�Q�Dl�۟U�b���U&�]�s(?o�QP�`��_}�����ZC���J�-Q��G�K@�k���VAZ&H����_�A�ʟLIW?��l�ꡊ,�M;F���Һ�K��K���@���r�/���\#-T�L�㱳Ϸ�A���$���O]?TM��]�fS�BE ~Ɯ����}F��CW��~��1�g�1�@@ޖ����u2��R��P/2��a	)�
{��U롗9��e����"�'�
�f�hvԸ�0����2hE�����z qc{�n!tKf0���*���y	v���7L^q��)�5L�A����;|晽�:�9��g'��@���(*��Rp,�2��'	@w�h�S�W��_��ê5!Ut��&:�Z�(�Ҟ�k闩������R�RL(�w��1��<���38.��*�b�C�*
f�ʄ޴��c�7_R�k���b�u�]�	��=��������p;^vh�m��Q��W�` �O`�����Ǥ�?U�+�W���̼.�ᔎ���ŷ*�:V��J�B�7
܌7��i���!02V�x�j���'y[�N�ؼ�jh	�D������� $��e�8^��@Dl�&��i8��̱�F�<�*n��<�B�9ڳ�L�`		O@���H�H�}����ʲ/(�^:f9��Y��	!�p�vD7�;6�ˆ�zHf'|�:�%�SZǏ�i:G��8���]�5H�-��]�7(��n 	c�$��ދ�����ӝ�Ѿ��#��_=����]�����F�hl�=�7_�	��R��ǟVpˆ3���[��'������FJ����/�:���q􎟿0��g��u�r2� ��*��	���l:	��h~�$�ўJ��S��(�F�!��Z'F�EP�wW�|�(<��Ӛ�k-8�tJV���R�d�S&G������I�{"l��fš�2��t?:-(�"�q]��<��2���d���H�(L�7�d�0��gT�����:�Ae����4�ؿ��M��@?@�y�.mM
&�����(�&>����$��(�I�b��������z����z���@v`�ڞ�i�ɳ9ܚX<��x/|U���rS�������I@��x�����}�G���7|�<šڳ�꺯��[�೥q:a�"o:�p����r̎�Pp�#-X΍<�����*���OjJ��L�Hf��������Љ��cI��MQ��$?�B�3j���m�TQ�#����;�-~:�³<O/���S.v�.���R�;�Ќ钦 "����e8�~R�97AM��� �`�WX �ݴo�aM����JX	ٌ$�3y�<?��FU�z֌*Ml�e�H�c<�!�&�_h�}ٵh��41�]��V-@�`-;�����Cn :c_�
w#6-ӝ�D5�!��8%�����aM�0�u���*h��{@8`���j��R�Ͷb��T�Wևs$�Y5�'8�
-�dF*F�4�ģ� G��+��t�4d��N9�i���1��-���XT�'�`�{fp#&H��ks���Θ�r�-������({T����8�Z�9���U}bb�`̕)��g�,7�	�_|B��Œ]j<oaDl��Q�F[�x7��k`�j����<�SM�y�g��A�!9��P�)���+���ŉ�89w�`���u�:Ø�O�{=����3H�&���o�Z���rT�U��=ҹ�	\&E�CU��u�����U��b�����E,$JnX��m�����m��|up�R��%�K���uǂ7���@�(���ڑfH P6΍�G~�����C6~�f� ���43vv*�9V��_l'�����Gi�'1NV��3׫bJ��J��Hg�uL�m,�ф�@�(���gQh�uVJ�-=�������]�e�\���P�E]v4�
ՊQ�V�P�����%_�1��@�s͖�*�Zv�l���݅�3#�x��:F�bi��$�hC�H���Ս�v�5�|�޽��0���!7m�:�6��N�A���Տ�J#D�keg�x�;ZWzSi�n��{˞C�(�PS�0��Dـ�zZ�H^��o~Vس���.[�R�.g�E����4 ����T�)������J��lX�M>�=��vLY�%;Ģ -���g*��z2�O�~�*�%�o���0��������!4	�w�(G�7���������R�ߵʡ�9�w�&�m�vg�Z�96v�
a�=�$q +m��g��r�Q]V�\|�S�v*������1��5v�=U�g_��;�X{Js���7��|Wۀ��$���߅���K�N���ǗS7�?k�����,��pu��k�r<2�G����*�l5��K�J�AD#�T�V0�b�*�
��m�u��������3W�"�����Ƨ�M�b�u�Q{�cC`x��+c������+{�kدU�0 �S��A����	 ����J�{���^��6Ђ��,�����,x�|!d0;��J�N:O���߄6H���Z�&��A��p֧�:;�f��
��΀�C��v~)���F�I�a����,Woxb1E?��ξ�[RRԁ��;�ɭ���V)���Ω�y�B��@��s�_TծW��u�"�@�-��{�2p�-U�r�D=�;}7�cgX�/����g�W�l� )�OHi���z8%��(3�`��r)e����R/}�+���D�J��� ��gqk:C.ⴀ�W\��5�7����C�~^�O\�v�IFcACՆp8k|�_>TL�i�d���'\�ı�2�7�L��e���2��"ͿM�b#af�r�s�s�QE:R����*#�rK��EZ������c��׫��M�P����*"�08�	#;w�V����G_��"���`.�U-�=SN�x�{�ԭڳέ�P�|e��h�%G��))�2��j�:�.`���)�K�G��}�(3>�z��Ż�תh�c�.�q�m!l�yB�CrD���n�e��8`��=J�xxѶ�r�&�wy��:Ƞe�X�/�O�piD����X�:%Kg�,<J�}B��4c+�i{ϵ���9�gPf��ї��6������*8��M���'"�o��@O/�A�R�0�/%�uC4뀫��d`�W+�}n��~�}�u�r���K�i%R�Rŕ��A��n{i�sI�c�A3'@�+*b��~��l�#���#6�/�����63�U�S"�<�H�,����>��S��l���/<�l��.�.�3I��T���s9r�ei��[�����5܊r]Xԑ	�B�zw�ƛr��i@,ɢ���,r�H�e�:@s�.X��ηL��/�}�3d$����}r����cEE\2��
�_i��O����oX+�f~��n���:�T�j5�D��cZ��wt��{0����̑�ҽ�5nK@�һ��F��O�f�S�c������`���_�]����YI�@��jiBg'`��xF����˲q��w�W�"Og=����.��.{|���
�9p^�ĕ>����W�DOf7e�.�-��Ѭ�^���V��F�r>=�
|ja�"a�vV|��Η�MG����,{�L��ɝ������q�@b�DdX �%�o�����ٮ�#��.d��/��'� O~���l��o����Y:J�$��|���$`����^u乴�4Q�� �5�L5�b�]x���i���X�-4����b�b�
M�|IxB��n�Drzv]��	ԝ�⬢�W��TUVW0]�1�i)��/w���&z��~��uT�1/|��ݚZ1,^���cz�8�vv+[sm?asQ��&��vqnD�� �
��+���^����sV�Dj?m�x�K�X���ҥ��F�w�-p��0IL��P3���3�T���	N]�-�Q-i�X��{OA�+��	�8�T�u�l�U�׭-�9YctO������, ��y�zqnb��Xڟr�&�S�@Xw�!`�b4U^ �\?�����I�'�;�8������u)�X])&�Cf�'"O�<��I�=1ᢒ��O�39}��P��1�4���v(�
��c	R�a�U(�v��o���N�xi-}y6��6~T��+!$�ً�����۪~΃���?֨�������ˤ�r�!8f�}�)u}����d� ��%L��2s}}x�V�s4*}:�\����8)v��t<�2A���F6�n���{�X_E�'D~�����	w�^:*x�&
���r� ��	�Ӛ����u��w�����������>Т��
7m��vll�i�D�tc�El�k�fAm��e).�3�t2�A��Y"�ʢ�s�g1�]>>'�񁂤�ôod�pM���jT<��@�D��?�|!�6�ZG|��uD!����&~56ygmXQ�7
��*
��]�v�|���Ťd�[�+r�u�� �m��L[��� �t�<�b��Acu��"Dfr얿#e���������S�t-�n��sax�F���x#F��{,��L���{�?�4hc ���S  ��/�
w�����78�`Y��}-ߠ>�_лg"���Dާ�ȍ��0A��8�,��O��
A�sw���A�*��J�~퇳 �,8�V:��*����C�JW�A6�t�v8ͳ���d�G33��΄����q�ٓ\�Q��Zc�,������*�l�,O�z^�pk��9�� ���B��5p��q	+ 瞗�wS=�B��\U����U�Iw.�$6�n���.I$'�DP$���uŜ�)̬ɤ<������ѿ�*�o>��������U�yo%�-Q�'����e2ٻ�+2*V{���M'�!'�x;��F{�|R��w<h��x�v~�	{C�>}�>�M���d� r�����K��L�uX���2Ņ��Fgv�� �Y q�����c�mz�Ȳkg���	�łO��#Y�z]���t7�E����R�5���] �QK8����<,s�����隭�4��Ͼ��W�D"%�A��T�ҿ��ݮ�h���$�|��D����R9=~�fn�#0C���a=A-,&�n�Z�=Ĕ$r�q�
-y��|���r��������X�Ț�3G��e�.�p��o��=����1a�T˾���Gka}JP&�$��O����U��6����_�h�poc�����ū��O%yW�O��3Ze�H/I]wB���;"�étt���#RM8+����Ž?gٿ��3�[߆6a
�X$��{r3_2�w�p�����<3�c;�'
���Μ�9�]�U����U�V��iI�G�d-����:S�)s����>T��'�5_�iI�F)�Y�F�o�� H�����%����"��^81�f�y�\�<���(�a�;�P3֧�>O�FI0tk�#����Pyt7�O��ڰ�Y�Ѷk0 ����q '�)[��Jz��*�0�m4��&Bm4�֠�@R�6q[S�w�B��$��*
�hyrq�4��՘
��(e���X��Y֡�Ӹ�!(�h\V� i�ӂ��7���xy@{���d�ٺ���θ@:�Iii$��W��K[��4�淲s46�!-5�>��O+�̰Rա�3�W��'ǚ�2D����:����e��w�B\�=Ӹ�tm��԰<�3�x�[���8�asl�
G& ���)�2�a���$Q�n����h�X�kx=�~��0���O���fҚ6�/���"��' �ʑ�y�z8�Vf��-�	i�-�4� 9}X�2"0���+ۂft2�]�}>)Ѯ*�+�6��<'rn�9�t�θ��߽l�i�3���o4��!�Y���u�����*�ۤ5�tH�AՆ
�.�h(�풲��F������p\���Cxm܍�-���]P7���	3�:�gSwVq��W������4I0�Y�0��[���[�h"<\�7j�_��(�}1��v��a�:�}�������6B�������=ʳ��\|�^K;��+Ƴ��.K
��]X��\g�6�P��˷V^;hDCݜY� v��m׆p���\:k
���Z��֥���JI���DHJ1�?V��JJ��OQ5/��6�g2Gb�����Fxǣ/��Q'@q�Z��[OP#��U�s-��)�
Q�J�iZ�Y���4��.C�g:/S[�@��ϊ�xor�������j���ѡosL�4��+1���It��ӝ�1��q�i�X/bm���6쁝��\3L�ܨ!�F��X��z��bD�h%�	č&����� ��v�iJ�,���}>3�	VO�����5(�:w�S����L/a*F�ͳy�ڝ6������G�j��g^=UB�B8jz��W���K��4�$�d���KJ ��D�Ӿ$]4����Z�Y����|u��7ۖB
PH&� �'5�Υ�ɛ(&�ae��� #L�����6�����#�[kr���P��8R�wD9�b���F���&oS�� 4u��I���IwN�6rמc�#MD�gC�|��V�� M�q��*R�;���:1f,�PR ��Ƥ�I8���(F?���I�a^�Ζ�տ�X;���}sT|�6�hg��,g�Y�OPi��Pd�x�x�3��1�Y̳��wٞ��0-���Q�n��h���P��C�7p�L=r���>����ڸ���E��f����b���c=P�Z@ê����2k7"���-�$�x��[��5�k��}�?��u�D�JW�%0�ɱ�h��ˇ�qP!/��k������ &�*��E7'�ؿ2��<jhu� ˝��!��{.�5;�Uq[�����.��[_R�A�0o
�U�sT}��u`F�
-������ߑBto Լ������՝b�/\��w��8��9��إ��i�����v-�K2�fF?�i�Ta��4Z����`��ޤd��#`�R)�����IX�c  �� zǐ!�:[0^����>M�Io4[�?l�N�ӿ�Qt��3�H����������~i� �N�
䃠��� `^n�zm2|Y�#�\��L��M�I��e��$(ft����\?�LI�+��K�F��|2��+@�&]U�n�,��+�8\���A��\>�]a��h>\Z�8�l2F�ed_�z��"�T�_��i���s�z�Ur�bro�j\��~e��h6���Z� b��\_݈�l�m��γU���A������������ ���t<&�`G}�Ӊ!�zz���,�������1[V��G%)9 �/I)5�IcS2� ��wے�hY�N��6�C�mkG�1���X�.�C�"�
+��R�66�e��L�<�T�����D���0��]#�lт ��I���������l:˞�/.�����=��B����t�T���Um�g�~������w����Q}
��4 ���/)P��ћ[Q��}@1�q�9��a���✠"MEc�r1CM�W6ϡ������)O�T�]=l�!r3�B��^8ڭW:�@�����N�L#��xfsMeFD�e�3,�4��]�@��mM�MV]'��������I�,�"h<\�q�H��VwFy�tdhQ��8�L[�:[<:K5j�?2m�XP��9% ������s�J��2[�����#�wnla8cc\�y�&�� ����;�dj�N)$*5�!}p�p�я����Y+Ƅ�k�	![�ڳ<,��c�;J�f��U�l�Ǉ��/�	�W��W��(��7f'��x,]䗜Ө�Ō-2k��D����Kj��~��0�Zx���	���-p���x<�x���]%'�j���D7���Gh��+�C���`����A�1YWcP�k��*�]i]�r;'X�w�5�rQe�i�cH-Y�{t��^��<fw�����nw�מ���k&qSȑ:�60|�����?�q�yRyD��%�g��~����Q;D3u�4��az��#-!wD�_�:(2<5�V�X�4��*��a��Y�&��W��z��7��sXb�M���kX�����a=��[�^�n��pO�}Tv�+N	ɋ!|'�I�	-%���hQ�_mw@����&m�φ���5�1��n�ےzO6�MiA�:��q�/�3�z��k5�i��ϊz���y9�29Jc���MF���#!I%��6�?t+Qa)��\q><'于�n:��~�M�_���e�5K�z4	5Z+���[�T##���0��O��m���X��#���^{�9f��P����k�k�ߑ���R�/5/i���;��N>;m�b�7Zi�>$>�7����2�~{̚K�����[e>F�5�^󃅍R	��`�mce�w����������5�N+#7	��Ue��E2PΨ�Ě��GC���w���'��0O�����6U��%=�^R6�C�(%�k�u�MJ_E64h�0�F���T0b,pL�ye��������NB)ϙyi�Y������E*�><�^�(l 1?>C5���8�v�67�;�����lm��Y� v��F5Ճ�ך���/�-8;��۱�h�Ͼ2"^D��dyf���G�1k�"?���q�������i��.�rW���ŋ������i�!6�<7�C�����̋�T?��;��L��q+r)VXSm�ji��CA,˅nL���h��,r*����o���W1�%���՜w{�kp���3����kN�ݩ\���o�.��?D��<�D��Ȉ��t엮�#�;��2��("�������IE9�6��bxuɟ̗��V�DK�V��4��;%7����&���Ɠ<���䈧���ރ(�6��v)�z��;Z2�'h���U�V�=�P��Y�4���#�JJ��WM{ٍ4݁JI�>1��߅C k:/>"=U/���U"e] H�T�60�9�ʼ�������X�	�n���6����R����i�[�dV8��,le'����O&�u��C���⾤���T���oK�	��z$�D�Cxb���7�z� �]��1	�&p��-#zA���,��V�� �h���g�e��q
1����^j��!]MCxB�3��ղ1�%.�aN?~��(�tki{'���h�H
a�.��s�q���V��n{����j��|'W��1#G9X�Z�_"�pg�.����G�a,��y�|L��j4G|̠B�Q�j���$����(O�i6_7L.xߊ?v�����ȏzl�3O�%G�bk�lp��׈����x�?�8�sy�\]�6o_A��7�*O�9OJ��Ԇ��J��IQ���`b��Q٦雖q)V����|;�EF3I,��)�y}�THp�e�:I3 l�z�(�?7C�x!*��̷�j�54~D8��'�һ��0�^;Z# ���� q�N{|��v[�}�k�0��
ݞ���x�6��5!�
?�Z࠳9"���
	!�l@��T����᭯'�r>w�8��t�ę�/HK���E�jiP���  ����yZ=q���mϣmP�?9p��Kư-�������hW&x�/��é(E[c�1]L�S�!�K|t6���{�+]2�Y�Պ�ܾ��D�НL��!�ICJ� v�=o���R����P�g�ϭ�[�Za	�!��x�ɔ�� 0��_��!j��w����$��-���GȺdű���,3m2����gv�,8�!q���2�L^ĳ�a���3W�yvd���ƾ�2�ι���(w�j�`�ؚ`�F=8��P.2X��l��o�y��vR�C�`lo7<����G�P�p�z#�w���ø�th���Z��fo�i�	�Nd#�6�t��{���2a���a#���4������t�=6L20 �a���mc���O8��q�Mu�A!� \�N>��V
6M�s�#�wTS�(���ey�����1|�_�m^&�ze��uy��Ɇ���<�L`��,���}�G����I�*��Y��<�MQ�tEB0�m����S
�M�?��h`;���=�+��:��/y����Z(Xr�t�Glރ~l�-h���Rat�`��%^*�Ճ�4��v�_����/5����"���28�}�?���4;\�p��
�����2[�$���y����N��1$m��si/.�O2ڸ�d�@h+[YZ�q�w��X���ې'�A��ە�k٤�{���;�P���Z3�5�HR��W��ƣ����k=06mLMa�~h"���p�Y�dL�}��I��D����v�E&P�o����&,�2�L҆o?�ƞ��c��j+�E"4�Ñ���&�7�"���W=��Z�N���U��0�l�8!��VEiY}:���G��
�ٟp��l~�H�D�|�S����ۋ���"7�"�+������5��k&�nAEĔ	�fk��u#t+3���bK�h�\1���i��ҋG.�#�qbg��"����`_�?^�&_� �yGARƥ�I��+jj��SJK��	3ǚ9�r��7t{�����=�O@W���@3�u�|���=JA�ީ�"�4bz�*N�.���%\Kfj��d-*F�сľ��*.��e͖a�M�WC��k���g�(w�� 
x�+�C���j)��i�l��w�Y���t��p�S�[�wK����r�����A}	��(�1��LC��$�d׾�B��-.��b"��껴��]�/���օ���\,*�]��C��T���a�W�y���v$S���s�������9H�Z=?�0��`&3�U*?ï�`�^ �n�¼�)N�>�ׄHԠ8ܼ����c�9[����4ZL�Y��GȈT�,�Jы'AAۡ�����d�So���f�����{���-g)ME���| ��O9ev�[��4i�Y�ޏ¶k MgM2�m�b~��<T��~�L�*j����t���d��B���3 z"�
_���@CoXGZH��Z�P����ҙ�L�l���� �O�����E'�m�'�U�����q起�+�޴vc�=K�=�Qi�_�Џ�|���|g�xD;ܛ>�S��W9e��P�aJ���]�?\���������9O;_��#������/*��c�'���P��ϜM��)�˞{�u�ϧ?���	�~�XY�������>��XԀl�Ӓ����B�QŃ�\%;;+���x��(�m���������\D�i����v+O�;������>�������Ь���et��gu����`�g�"���<�;�@`-��� /�4������a.&�I��OUa��Xp��X�1E���+.Z�V�If���O�K��R���� �;-�9Q���{�:��S���%|s��{�#^�ĵl��5?R�S���yK�t��YM��kI��?V�,��� *�8�!Qԡ�����U؜���뷽�(�55D����p�B��	EC�q_OE:J�F3g��l���O+����Ov���q��JiH�4�a��5�e�Q���;�3������8�����Xp����4%wz�@�EM!_��}�K�n"[��Uvv	�F�-i|�#�iuv-|5��g��'�*K�;C�����#u�"��v��hQ��΢� Gb����p|�>�wc�M��w���Z��ʖ߻5�4A;�~v��ʯ1�?�6!?�2�3GEP>?��N�C�rpQv�A���'N�����T	J�
��W�!�7q7%5`�4vcAj�ȁ:p�<�=�d~J�h@�νTK�X��Tb~`�'�n�>`D�5`1��}�oĺ,�Oc0�# q��s�ϭ���c.\F*ΐP1�q,�O4'y��v���ʰ�A�~r���l^X<��#����t���<7��~���F���m�f��Ȋ����<���*9/\�U��s��W�L#E��<�j �V2��O��f%��?z�������]g��OD+���8�z�������Gi�l��-�����\��J�n�v�(>��⽒z`"A}��K�0k��m�h���τ�������͈U=�~�p�������p�h�|ġ�$x�º��J'I�9)q�g��z 	��9�D&&��]�-3I�!컍��1o�t9����>�]c>.�s\D~衣���.q� �d�Xf�e�����nQa�*/�j�i&����������g_��%��_5�3��wt�"#8�K�~�L<���0I��S��%f�f�Nw2d���pȋ�l �9V��Wx|��{U���(��j%SM��2��\��Ǒ�,7�M��>;z��ur���7�vnG)�v�H��Z���v�ۭ�t5ihv(S6�g>�*��X���x�(f>!�������Et�|'X�@�w���ݸk�45��	�HC�+�$�N��]~��?J�0ӄ�=�v
mM7��p��4s��E��� �ۭ�
�1w�U��(ڎ8F�JI�{�j�Ԟ����k��2��vc�����ƞ��\�����$�Iщ9��:���j�aF�u��+�=� �u�
:볡'�]��}y��$�UR�	 ��P��l���╈�a�Y:B*��\���N~җ�׳��v��WM��&n✜�{��[���
�4����r{}RM0��	?��ـ���/�$�D
�=C�h'oZtE`ikl���Z?c}a�ds��.~^���i[�b�M0�1.�xj�&z�Jt>�������m.Q&���w�t�C��6r�H)�lA�h�e���O/��pv�B��i���c�+2���#?�lX����P�U�e�ֽ�_p��������u� p����ռ���Q`�~�RZ�5��nc�; �R�}x��\`t����;�-2����sp��Q!RR��{�\�.J�'Ϥף�?��Z�,�cl��z�U�֎� G_��!wK�P+[?uǶO�=mѫ9b�?#�4:�9D��[!� %���#�� '��u�u��{�x�X-o;����*V��=���` ������:�Dҷ�Z���Z̦��Pqd�V�ʷ��-�􌠣�O���M�o�M�F�@�6��9�e��T��0?�[���'�[��"xRb�sbL%?�6�XSN=3�̤�(�rZ�AoW��zp�<R��]Ԏ}?�o�Q���f`��]��A�X��y��^�����gT'�,���i-��G�F��|��y&T[����A"���-/ ͬR G|^K\�}���	6�xH�P���S��(4��oķS�jZ��N�W!����)D_��x]q&*��K��*�%�Pߖf�#&��uE�����>�[�j%N��<#9���+΅]\H��=������ˎƔ�U�ij35�	t�܌��}��'��ŋ�G�H�Ah�R�إ���kCn�K�j(5�|��@é���Z���%d0��Ϥ�t�z0[����9k@߹�8�4̑,N��ٶ�٫��b�e�uYZ���<QMS�`:�6�w2��a��N���%�M&,��;lmm0�x�n��c��YH�۱�aY0���~�Nm�%!�'"1|#���HP����-:��@{k��Y��s��*�h��3 [�<���C#�8�ٟ��q�� Ґ?�]Bo��
�[C�R5��x
�N�S�hJ��K��Q�ϸ4g�/�xށ�2)�R��������!������#�����u#�W�4$O�.x����}mu��x��y�(�W:�����`��a����+�<X��ץ3�}�/g0nJNk�bj�a
�<��xO�$�3�a�Np�F��Ku��҆Ul���?��?�c���b$���A���qÖЖ�0�].T����F�ܨ?{�f#>�9F~�@�ɩ�W�"���z�E�D��[��zu�<w�a0�J��0�1��_%fK^N�T��p��'�pצ=���|Ή�Q�Đ12����O�{3R\+k �"wq�{/m����(���^`+���{���D�Al��O%�K�	�5��ߢ71���*u�9S
U�"�&�H���9�"!V	n��o� ���n�t.}��`.���?�)zS%�|ʻ�K̲ߴmPy��a��r.:]�{�8�sap��̽**�:i_h���1+vCPn�0ui4
@?��)��o��*�@c�z�)ʃ��v*	�iɬN�f�IE�<�dy�O63��)��Vܻ���N/_p1/��E�y�$1n��Q� �8�_�1x��G[��{*\x%mnRj�hRG|�_:Ha����ݿr�Tj�i'p.+�{���]i�^rE�B�ޑ�?67�r��r����6��%���$u�+�P��)��ř�H��	���U����3�I�uS����|*�<���+Eh�H�g��Myթ��T��	��,c����?�CzL��әd���8���п�i@b����@_�"U�ƕ�2�_��Q�S���{�_�����m~wX��y���K�ӑj�O=�'z��͍Ce�4�ɊB�	 ��d޼���2�� ��o�;J�;� �D4餕t'Y���l����"����}��Q;l���%6�ꦈ@d����7�
�tM~�L̏}-���;�.��[���D���Ct�p'�.��,a����F0���t�5�~�WУ��+�=��mE����\����s&ps�XE��,��1�NY���G@��������'H<6���M��K�ҽ�z�.��mDhd��s;��,�5�! @x �5�[;$fM��M� ΁6@3TC��bD̐N���0���*.�?�"<�Ft���Ƭ�0c�Q����~% ]��Gt�����*�]t<�=J�+O�>�@�&(EG�;�6#�^��E-����-$˒H���VcM) ���S��lw{�R�~{䤎c����=�=|F�ZY��������`E��{d*�g�����/
��  �� ��δ��$t<�]5l^铃�D�a��ъ��r*�C?ڂyc��Oa����"�<����A���'	[p����2?n�C~ ;�rS#@����b]��˻���d��v�>\2	}h�݇(/����S�����W/	 ���a��LDj��]��j�k$Qtc�u�C4J�}�'�����,�S���{ރ���1���.z��&m�еa
~o��׸���i�fY���BHk2���B[1�[*�+�����|��{��襨�{�X 0�H��	���g�_�E�o8�o�s��M��C�c1����hؔ��`S��7� J4�u؊�1�uw�JψE���a�ֈ�.����RQ�hpAF���0�i�1���8�4��~Ȓxk��Y��$��\7p�n�9c�4��_`� �ڱڀ&A@7N�W��(!�Э&��<������ն�zM�Tbz��|��0(��r�ӑ�w���`�i��C{"�XmLg�?�L�=kg/T\�f|��XyI�cpSt����q���īٵ/U��z?'������/Γ�_ �\7ܻ����R��n�ߟ�����e�m�gÃ���3��Y��սC�����8[����6���ٝw<��Δ.ְՆ������Qg�Bj���P���D�UL�rYR��h��Ζ�ӝ�V�22��22ޣ�G���_�]�9N�C�����5{�qNU���ʒ�1r�>!��Fc�*��{?{O�����KIS��b�G�1l
A�%�x|#Yy��p�-X�R��.�w�w@��s�>3�e�'� �v�|:wڟ<��!�A�I��ʒ��	��Ve4\��2�弄m���3�7�3f;��hk���fj.`������w�ю�{G�m%�`O�0e��CF˃%�Z���
��2@�V��b�/�l�7��o������3�\e�Jó�d�6��F� a�G^��2D@�a��Ƚ]]�:�A:�q����gE� �I�&LH�l�����S��;�!p�w����1�Z�Z��#-!��R��}x`(�ғ<��X��w �VЙ}Z?�^�9�E��uR�԰V��K�t��F���T��!��L���{o�������T݊�	��-��0s[��.��ok����[)�)j�k�'o][�S�t�4|�:���P�';&���Z����<�)���x�c�vjҞ��c�9�+����\�mB%���F�HW���oM�R-i_�=k��I�i��ײ���B���nEc�)��`�\#_���
N�-* @%��� F>vp�}���~�@��al�Ǻ�ںcX܏�4=�����$~��G���cF�	p�d�d7�<K��6Kd�'���̶`���(A�]�%;�
���.�i���Nwܥ�_�-A�6�]���Uc�����haě�4�_i/��o��_�`�@Ԅ��f�"W�xss!�Ů�͠�Ja�8Tt��E7d�i������Jl�v`���;������������f0���L�<<n{�}��p�#�?L}O�~.�]+x!B�j%��������[[�Jk��8�6lu��*�%�3�{�+yJ	��*4F9�㳔��F���b�Vn��6f@�z��z���g�EE�=�H�%���#�/����.��2�'#li�u?���iM�i+���4]�)ʩa^�	�B-����#��n���^H�
�Z��? z���Xm���0�b�5c�7*�6F.X���.���/B�P�*b�����aE�vF��-n/�[H��6���J%�60��"7�dl��Cϼ��.SG96;X��ŀ�+��y���-�b�t/V%�(:=�5�3�<�x���) �h��0�����8J��<t�0*��
R��3�@q����/���8���i�g4ꔈ�%.�5k�u	�}N�$Rid>C����w)\F�Yo$6� ��h�������`���_�|�s�B4�*։�����J��H�L`g/��CH�*��8���N�K�����'y�AY�ר]ZiUYJ->9XC�~ ���!܋�\��r5�u�� X1�m�ƌK��	KA4��d��$0�'�aA��^7h1@�_�mu'�Ʀ�u'zA���I�(�Ϩ���F���2���/L�&�z0�$8yWU�hV���Bl{��^� ��o�"E�����;Y�_�^����3��(��`͚ �,�h�K�7�͌ژ�����N�+�$�PT~%���{�}:��|~�M����嬚�
MM�z�O�SOI�p�	�z�J��H7��v˃�w�F�ڳ#��Dʪ��*�v6Pq��ϡu�7X�����3�,._?i��#��	����K��[`VDf��rD������im�!^���o�O:�1��X1@��Cn����x�v��\�Y<|����Q�톶8��۾�T��P���"K�&����o:�h[���c���������A�K8��&S��fQ�pw��E��;���L�M\�_P���H�yT���Sd1��Wo����Y,-Lw�x0!ٛ�Z�)Ět�JLy �\P���^�y�h7�s �3�p�!����o�`�����y	��#�3^�0eRb��Q��ht�]һ�/v��)�f������
V�������
�z�I�HX�x��٦J�ڒ/�f�OGw}Y0g�줷���^��%��HD�W���J�Y	��"�9�����*?Ti��a��-N�b��߷[Kt�wĮ�ɑ5����ft+ bQ[^\�����#��]�O���neKƦ��0��Zu�2T���Tto����Q��d�m��6���w�JC�A|���,Qj�2�5����"\Y��=�3�އ�O9�B%M�Mꄕp��]����C���#!�G_x2!.L�|<{K�k��옜l^ۏ��C��������@T�����䁇D����p�C����Å��}�'���mP�3�З�����uVFL)2��|Յu3���8G�A� ~Jl]DOn�!2���r��5�]�\}-Y�kӔ���H�V'�}����7�n�jzdӮG��Ƕ�V�F������~��H�����Dv&l*���A����p�75C�/ײ���tV:n��I����G��|�)�&%��شl]-�����ג�+��3��ɀ؆g��i�l-�ۻ֒NѲSJ����ʮo�"f����,�O�CU�q��R��%sfİ�n=I�����J�9t;��&ƨ��Ed�y���-����4cGHl��<X^�N�6����Ki|�+ž����ߏ��W��!Θ+�+�ô1��Q��GSՀ�������xR7���~K}M��:�;��]b
�XV�w����׸�pv��Pۋ�r��y#�?�?|?��W����ڕ���q+ՙ1?��Ƿ�")2h��¨(����v��4����;��&]�>n������5s"~�k����e>��K
��Q�3��2iz�jw��0��沅�/���O�L��NT��&7�2�M�	;D��>�S�c�7'b$�V,�#ɠ����fɄ$�5�#֒�9��^����PF��8��h�E��#�}����ATY�3�������G_D���!�ͨΫk�{�紀���v)e���&�,��v��b�#䂐�"s�An���Мp���]fiT,���I�l�}���/��#&���X�S4׀�\�I�z���[V�E��8��>n��sɄ~͘�۵O�f�e/k��`q�#w�"��1ֆ!�(�ĝ�d\��9h)^X)��u<~�����o!M[`��[�5��f�;�,�����x�Xb[�Mܗ�S'ٴ�ik��l��X��]'ʹ��}?��������ɴ��d�_}���'���s�'=��9���3�:��m�w����^���w�%��c5c�	�C�`
%t�~W�n�5��f��j�Y'�/�8�b�[�X���D�B�Mϫ��a���"���aͻ�@�?=RbL,�.��
ښ����!�����z�Tu��[H�g������
�S*�2)��Q�&�*ZǪ�0\��0�{�#C�0�CDd��SZ��x`�b>d��t��S:��l9D7�M�U�s����V	�lˢ
/�ɐ�}櫌~x���RgWUϧ���mٛ����팱Ä� �"o���	�#�x��1�Q�.-%��}��5�I[Y�t8e�ī��L$eKTJ��ު�,X!�E�j'M#ug]�oڷ`���u�Ǣ��Q)�ǲ�n���f�)V�0�ɿ1߀�������Y �tO��T&P��֠;�N�����>w2a���Ñk�t�w�|�qĻ߅�D���V�ቼ�[�Y�4��$��\6Cd�_Q�iBnK�K/gaRF���dTi��*���˔-���fk}C�@��X0��0��}��d��"O
kto�g�B?ke���Qw���u���}��Fb��e�,�Z+_�,�A�hXI�w_��}U����|?v���|�UXSV�g��n�����d�����'�����n�M܊b
=�}�!��zٽ�a��  A.)�|��lc<��U���9����=�q<��˾�I~;ſ޷�K��G��?">�����t�7N��S^��j�~;��Ty	��6ݲ馼��h�6MȤ�	��;�.�Zjh�����{%V?�98L���">e;��S�˳Wf�4j̉�l�y1�V"�,�r�c�8����!I? ��K�kW* Cm5u�L��s�h��M���Y��B*�P�(WO�S������'a��Z��U�oV��{������98a�+�݋��Oj!�ɫ<4>��8��f-��^`yv8 \�'SX���]S�}ҟ�w�������^d���slHw��:T��n�'�L�Ϭ�r��kF�"��B/�해�Qj�d�pY��V$j��#ϖ�ʡ���[:�F��or��pRt�����z�Zh�;�!:]�f�}pk��5�����T�)MdS�o��q�j~� ����O�|)С�}}Tgj)���C� �O�ߜ�M��ҫ�^M=����.���)Y�Z�IX,��7r>��kƭ�GUw�"�nK�{V-u���:\K,�.	��@��9�c���ٌ���k%�d�����ti�K�*��M��<~��񁮟P!գ2�+*� P)���l�m�U=�\-PQ��&i=���׎��9��7�(�8��/��Om��͵��R��}�8�cPO=�����&���PvW�m�}Is��s��G?�뫈��̎�I1�ڎ��q���a���Cc��B�^(|�|x�Y�]p�� b�cTL�Wuah��y���K�y��Au�g�����:!�;ɹ��B@@~�Y[�bӗ�����_���1�1(�`Ħp���g0�e���p�C.����>���M��h���`a�{���d�o)��k<͚���)}�V%��L��γ��۵iY��3��w���Uj����ɕc+iĽ3�d�w<`I��\�-���O+�+d�=���r�?W��U���<�8l��T\�0�t�o)�������	�v��Wk/u�5�����[d�|J�M:�+�������|,�}�o��������mu��Lp�!���b��J��6�d��}vY`)����>�
*�Ù�5��h��4%��jGқ��q[�5����5������Y���Fɮ����'I�Nc��hsŢY��uf�����3��NW���E���@���#��r\�C��7ª�--��=Ԃ�\�����'d~}�F-�r�ז��Q����m����DL}��Z$�4/��{K�Rd1$�u�a��Wh�G=��ew���qл_���4,@N2�c@�_ T�F�wO	�ȷ��2��� �ǓA����U�,��.��5����r)O^����t���M���q��ka�k�#��2�����RK�ͅO���g��jAnb����������`L�|~O�}!��]�p�\�<uo����֣�.�fl�Ju��y�>.r�/�_ڑ�6�Ki�7��F�8��T�D1{,I��:p�&����h��U�3SWZҖr^�`��������K�*O�b�ɨÖ>�ī��GP�c�ޮ�A���)!g�׊�-[��!b$��?��!׮���r����.���d���U��y�P!b�Rz+�lԝH
@�nk:��G�v��r��m�lx�|�+i��f��2'��H����1�DD�E�&��q�c±��C!<�X�|s4�Ψ�-YRP12Ă����Vu�_D�����QV�Հ�X����}m�]������tI�{:.JoV3sݪ�I��Z�}*�,W�e;�{�Ʃ��?%M8y�~�ٍB�&tp
4̃i?���Ö��Ώ�{>�FK�!��L�/:��7�vΘ�'H �k(���8`�h&�Z��e�
i%�}��b�����8���l%�q$rQT1Z_�������3�;q;�ӟ��������j��E9&X)�)
D�G�ߞ��@�j��C��Ls>P+HD��s�e+�mݒkp�%o�| ����D�,�k�U�,���u�5��D]y�n����D�c�p8�k��ʑ#\�:9yaG
.#�YK��~��9��x`��B Q�;9�1��;�q���������o&R�p�mU�* c�9y�-��Xѿ���Bg�:(Es����0
����U�l�� ew�I���8�Ф+W�!`9(j��f�*=���fGIiyVpL�uJ\%|A�㢣���������u
|!Sq�ؑ@���,��՘�_�P��,���h@9�	�)RH��p���:��&k��N��5����� �������w$O�	���R0�P$MY�p��)n�;@�!FR��Ajy tC��fV?O���u�I�J~�tP/��z�N�=@Ӟ�ȣ�	�����>�/�?cBZ6V�������h�@�7/̑��E�]8CL*梜{#���n��ω���
��:�bė����hR��w�Y���L�m�E��ڙ��D#+ٵ�����[���l���q�)��,mJM��� ��Z�\R��z[L6H'�y�ᯃ2�z`n}0��x�rz}by�V�g�����5qJ��p_�?��.".�p��rH���f1I���*XP6�ޢ��K9����3�0��t��k_�'~J���Gc5n�SR�y0̕Ek���d�E���{H*)_��n����2�Y�����W�F������P�X���Y)=L�肗�h�z��uh��ga��K���L�]$�;ȿ��-JT��>7��w�_����>��j�����-l���:/H5�k>R�=X�� /7�O�Ӂprϗ
���J�޼�z��Jt�|���u���P����%Űj�U����s#ɕ���s�s�c�j�
##n��ߴ229J�-�[V@�C�����Gm?����h9��յ|���q�	�T0P�G�	�/XRb��L���:��m`;���5�n��͂7�1^ ��K������r���(���jL�tv��i\�ȕ�Z����=�q�- �s�4�F�9|g���"̂��T
ħ�=��菷�d=Q ��j<'�?ʇ�I�z�.����N\��!����5�U��io&bm��p��`���iC�k�}�dW�B_3HfpW��u��u׎�5C����Jx1��b��/�eW�K�h<�(���,q�l�V�ܓ��������^��-[���D(%?3'V��~�q�ϳ���i��ǽ�%���">��3� P�P���x�"���gmQ���A}�����p٭P:~�:��OpB1j���'�#����q*�p)EKq�ӓ�0-bEy� �Y�;4&)��͝��V�k�!��62nS���b����9�")R;�J�0Ra��d�%��B=w��a}�B[T���y���܇����F�������1��e�sb��vO�pU:��@?�U�K�*���kˤ��7�wK�[�rU5c��r��b�]�V�nu:N���c�mn��l1m���:��|�Y��7]�oIp-�<�5�� �Aw������Y�\��-������C�03�h�O�(zc�ǉ�r7��a){+h��Yh5AP۹����7�H������DǗ�_�i�}O�8��F	�{�J��*^1�Ϥc<z�y����"?���CԤ8��`!�^Ҙ�2|%`��&pc#l��~s�G��w�п(��1b��-fM[����S2{IG���20�(��j�^�f>(�/�%��-a�i�h�ݷ���&B3��@&3�)^O-����ȜY{JT�:�~Rs��.G�wE�D��%!�-d����� tͣ?�F@���J�y��*�9��������3A��J�A�}�����_�9�L	_ޤ�-�Z��*,���Psw>ڰ9m0�ҩ�?�W��|�z�1Bi]�$��*���E��T�݂�`0�=���IuK���,���yꘒ����鴘�Q*�����y8���^�k�ě]�T���Ec����~f��HT�4��3��p��K}*��h�y���wHJ�hE�|����$�>5��\�VD&.L��7��$p00�u>TP�g,
Bs��p��ou1���lt��Y��*����;����6Ф���� ($}$�:�.[J@��x#�;�7�n��Y�B��҂K��K�:$��!�������~��x���W� �Q�w��RI��K�ls�[���J� zĈ���l�k8$@�N*���7µ�ΤT���B9d&���!,q�1� ������tZ帼����b��^�����EAK����װ� L�� �J�A_�6P6O�.1��L�=�{959�����:�������`yAp��@k��&�"���0�cC<���r(+)�\�Osv�Xf�hN�"��:e���:�*�Q�t#gBFj��P���/0�Ɔb���;ˀ6h�R~���Shb?��L���&�2��%888��$�����^0u�2`�ʋܡ)Z�2������\���� �6@#��	����d��W�V����qT	m�?��he�h��Uf���������t��>>�2av�����T�d97���4ɫ�YH��V*��?��0
NN񀆶H�l*���U�i���s��]� �ػK��|�LzR����U���^�xrXT��/�$�B�����,Ѐ$
Jj{��k8�:�&�J�NO�qm�Cw�=�۱N�6y��_��&!�$��ԍ��8�C3eLBn�'��!0W�8h�:1v�/�M����QE�I��2��ʢ{���:n���7�~&X��xAN{.��8�I�3f���[�L�e����)x�+>X.3� +,�,�Ҝ��(.�)�>��xrɈ%G��\�����?4F��>��t�#���#l=�{�W�gk��Ǝ �Qy{8]P�P��([��=f%&�6}�0�	0��4 &�<g)����G��O�#1댕��x�Q�]q��m�UbSq�2�L�"qm�6s��,� �QG���j���z�c�U����;\�j�(�~d�W0��;*��)'�F�E����v�XG�\�p��\��Ӻ�PD�تT���$H��1=�Bq���[�x�Ӓjр6n�[u\�<KZn��N ��\ҙ���|qo1_���\��(��6N˞+s~�-?�Ch���%csMZ����@Ҥ;�����y�r���l����Z��4��q�s	v����u��+y���D��{aw�c�	Bi��B��e�h�6w#9�憝I�8�
����(���qw�3��P��AǞ�������Z�W9���}5��o�w� ߱1����iȽ,�ܞ
3Ȃ`l�簒�|25kD��+ly�!��i|y��FkpQ���gRF�?��y����l�-E-o3�A\嗮^ \�&��A�j�B����8�32 ���錰ʓ��`�����	��g�\��J�S�����X�������僃9����-��E^�4׷	��䲇�E̘_p;��̿��(�8��C�G%+o<S�?j�M��H�{�SZj3���A���F���Li���9m�Ů0��Kl��ߣn*�J��� �jK�A�b��&ѽY�����z��x�Ɍ�\B� g"p`��AN�Y_�A�6��p���f"�J�(�i��q�*�]�\럛E ��ZvB�2Q�t%�}����~�;�o�'��"�����m�2
���=-��~p)b�]���1�����m�RΏIڞ@tc*����a�¤�86G>��&��}��$�9i����~�-_Ɣ��-n�f�-JS�X�;��͘G�&t�H˄�C��H����rh���)}���tSA[L)`	���}��\�"��L_��F��}�Pew2p�F�l�lq�u.p����ؕ�2��%�&Rʚ{���r}
�e�������C��%$�.�*�?%�6!Y-��r���4�n�u�톨�i���~?�$��}�9��=m�KBgu���h(�1���K�m!��Tfx#������E����Z&��,3��P ��}��,��d�!�8��Kv�}��<j	�H��օn88n�;�z4���"X�\Je:�9�:��j���sp�D�p�oV��+[��G�O���/m����R�^T\L�貸��ۄ����6�������������թ
�{�����L�F��D�f��ӿf��Ω�/BJ��to}2�j�s��A?���̰�̎���`sW�	x�� 7��>�����9�Ӄ���i� Ǜ�����釤k,�%�f^�����J���pSN�$	�*PQ#��c�F	�>�\i��q�+y��]��ns������4���Í��ޛ���c�Ս���a�?�H���-�0���4��a R�h	���\���Y.�H���q��,���f^�(Xޞ���|��Ѱ
���}�V��PC�"�ٽq%3����,i����@!mQ�SOo�ice���ҙsU��R�}������=}������zI��`s:O�5����Ȍ3Ǳ�qҶ[u��T\�jb�c/V=�'��Y&9]j��FI3Y�'�e��޻ 4\�����T�c�ň��_�C��uo���[T��7�9����*���!��z�Z�}G��Z�8;��ŭ���K�	B���e$��V��w�5��(c�S�`]�)��xR��J�̦(���-Z�2/�ݚ(g�����j����j��/��7O{X���"p�"�la���\RgS|��9��<�$�E�Ks�r�\��v�d٬w{�Չs�N���V��
(�C7z?���Њ�Ѽ���l�Jd"nє<MN`Cs�r_=��+�z�uYL��(�X�M�/7y^���Z�:�%B`���{�F�("�V��ϕ@�8����#�!X}�{p�݂%����ۤ%�Np����M{��K��c<����4UC��t�t�R;F���(Gu�ӻ�3!4��=Mdϋ���x�}���^ZN���GO"�g���1�܉���^YKC�W��Z������!&8$L9)6� ݮM^g���C$p�n�B���i^C��x��� �x8�ⷢ�3��A-q��{ t2����!��,�{Rq
`�ؐ�S�A����G�}^�b�r���� )��Q�"�t���2.�)y�a�	[<���$5x���n��0�N+)����f�`��䛽0����%Y��~�p�L�~��_Fdٞ��h��%�yHL��ՠ˷��3�U#��>�y���`qR/23�@����}kf�.�_�����5�"�B����3Ć�)�t��dv�V`26`��Vn�NE��^O�M�CVad��g߽���i��j�Nֽ>�qa�1����'�x|�[����Sl6o�J>����O����f/�gRq���hh���<�}T��h~�:���j����b�a�g�]/foNN����#S\�`}\s��}W*;�y^���D8�&%�T��:^ �;�8����C%��&λW$ݧ"�,�͈{�s��f�E��'�_�v�07���ix.�;ƶ�EpgrJ<�>w	(�ZԲ�Ɠ
�F1I�-*L���wZa�̚WF��!yCt{$g]ʮ䜺�Cd�	rð&��z�A	�������E��!uQ��>#�[E����])������z12D��w�*���RXK��֎W�%zw͍/i(�fE�LC���7��~��g���m��C=�O]�7���JWM��ju��:zNo������ƣ���uG��ԉ�zc9�g���l������h�o�����y�JB�(��1��m.��t��NC.ۗ�>�
xJ�������O���9�s��x�@Sm�$B(���2N�;��wN������\bj����c�&���,�H�j�t6�ߏ,�w���ER�ѷ@��F�)'M�f֦ҟr��++A/�l��1����jvq�P���<�7.�b�>Z��",�8Xu-iW�CH�$N��p����W�SKR 3�w	��\��kv��v�Q+�';aC�WA`H+�3�c' @�>�ar\=WF��t�׷un��!|X k6-��;L�#���̧򗗝��W�*K�;� 6t��-Q*Ҝ��6~���!H<>�MS=HKF͉P�N��v��TGܭ�e.7XjP�F���2:O���Wb"�wk���O0`0NE�l|̴�>s>�C5��C��Q��Y~/A�Z�q�0�BM�첦�`�_�8G���	/��2�=�zYZ ��h�M��8 �e�^ �OU�g����ZI�@�a�1��^~5��#@f5���U,��{Z����o\mn�`����ef^��W0���\򨓬���$�iե7�.���D�4��
�͆���L�\���[�֭���l�R��V@��S���L�Cj��d�0OF�lr	0;���]h:�85��R����vFR���|��	}6����&Z�'�^�S���:k�@J!��hY=��P��u<���Y��tD�[9/H��+��Ph��?�$L��~N�N5z�U��V1�T�ů)����\M�Y��4ڽd��*O��O��F- �XDŶ���x�8 �.wDVN�	���~L��4K��t�o7��@���E��U|�6�T6��d�qtf`(��(5/KG��ڐ� �	/�-j��vd�r���P]�,C���P^�ښ���D|2qq�D^Q�Ƨۻ�Ƴ��Z�wEN�9�zyX(������"/���PK���>̬�#�Z�I#��]�t�h�:��Q�y1G�Q���垩��_W?�)u|�7���B���k���U��7Rmq�<*x�h�~�7�����cr@`g��,Գ��f���Y�q?�B3�GK�A�.�R&?�1�M�B�ج��.��н�\��Hh��fcv[�D��!�zu�T
�SQ��؝6#�5.�Ƒ;�t�_�[^�ـFxgfu=A���>�6`�37{�� &��b�hxX�I�"�4و����t���X�����A큿�k��q�����X�XB�u,=HM�,�\�f[����h��}�r�wC�}�G���t-x�y���<�Q�%4��Z�˚���ۏ�gMr>A m����b��#�� �vPt8�8z�}�n���t��-�u�B�U,kƨ^�,�S�����ʽ�:���&r��,��L�zR��zĞ�v�Mq��JVV$�U/c�~K��D߁L~�y�6�*�z�(�:�bD���3�U:WmS����]�2Z8Y�)��'N A�:�R� ��N���D��p]`��	�<�H��'��g2q�l�RFߖ�����0a����������c�,���g,-z�}�8�z�I%{�3L�	�k�wĦ�urN�ɶ��%>��$K8u����?��]��@�8jr��'�����h�E�n⁉�nG�A��qf��=&Լ��p��mwF1 �%7� �f�qvU��.��Y�-�b�-IH{���{�����gU�Iay�r
��-�)��=�	���τ������� �߼�+�'s��)�U��p v�Up�R^V��x�RT�/��N[�i��`�?EߨK:a�X5e*�Ԥ�LӋ�z��yf&��:�~_K�"���'Tt�%p�5l��Tp�U��`��XM�/K��A7��!
��qμ|����a��m�iuY����ce��F�n/{YQ�k$��2*+^b SK���f(���.�8l��G���Je��+��C�B��m��h��0�k6'apf{Y}MyN;J {� �G�{Btm#
:�%B�#�Y�����Ɵ8r�K�3��	~����4����V��CR�R�뜒�4c�Z4Pn��[���ģI1V'^ums�
��W�?^`��.O>l��ي}���pR8<�|��c�����w]��2�,����"�K�S �shݤ�U꿛�OcK����������Aӕ��i�Ǹ}���l5碖S
`v��U��k{�M�z�"�늖HL*<�#m��Ws���IR �h�4<6�=�G�Ȳ�󗴱L�����,HuG��J�H'8�Z��{"��G��(�QJ:'�[H,��+q���*Uc�L��u3��OYx|]Y�ͫ���%ˁC�k���.��������W�O��.�74%�[�ۼS[�X���-��'IA�D�1�?0�K�.(�%F͸���j���B����G1Z�䪼�>��^�֍ r�rC{$�����k�X�\M;�{^��y	/�Y�e٨-�y�f�)rÞ]�2N'ͬ�u�q(��>�ȱ�����x�� VyOBtD�1(���?��X곊��:p��7}
�7���Ϫ����!K��Zi��F0��<,��UTB��R/�L��J���ѕ�f;�=�L��K2E���q�P�����y��<���1ץ�Կn��ęqs�D��=i��G����L���ג��M�!�k�Uze\�����<�%�6�W!D���)u<]X-�k����@3)�WQ�?(ෟS����[�ie;�2��H�q6��uL ��	'`��z�'!�\r]xȇ0�'P����7 =�|�%�O7�.P8P$�(�ܙ:^�A�P,�~C��r�Ϭ<�K��@a\6�R�J����H�Ьp��+��IҸ� I3�>fi�Z?����G\��H,ñ���:��Q�Ͷ��������%��F�ND�!r���(OMgv'ۄv����{��Y�J�ܩj�$ph���Ǳ_�_<e�[�[���˭��(�J�i����+��7�;��ay3(*��K٦�r��b�^���.Җ������B�V�0�\xzz�x��.^��#5�g8�˂"�F�.�ӯgE����Zq���
���[O3P�� ��u���70i[#)y�lS1-�
8�1�x�}Y��� �a�oI#�B�������ʆ����d1u�Y�S�~�˞RN�sb������\V�,h����a��|ixZ��N�2�ǹ���,�;���5�!UOii9�Bũj��:�e!���Ĝ�dP��l�	�o�j���Mc�^v�(>�?�v��S�
!�,�?�@w��wUCr��s�A,,�b���"\b��^��K8��B���rJ�@�dv�?��X��LADb�\�r'�������z{�ߒ2(ܦ�'���°��t�-6(c��g���w� 8��rbAt]z'r�5����NV��گ���f6�/}���H�ZS����]z��&8C�d�^&���V0��7!L�O�'98T�eK����o���T�Y��K�sǤ���>ϢrY��Q2�jt��S�,��y��h� ���������2س�O�䥟0�W=�{�p����7h���lN<^F�F���?<�E�V푩��(��y$/YM�i�f������4Y���;���1\-���� ����R�~���u�Q��s�S83rP��I!n:�ހqK`�|3�i��uYWgJ˰��!=�w@'}	�7q'ƻ\˗�#-��X����,8pR-��7���wߒ����l)�0z9��Y,-��oj�{Y�7�"h�t�}��0�N?<�Q���Yt8B|Cm��a�����"N��/3��9
�@��A��T��W�R�Q�<R�R�~�2��Wq<R9[٫�S8���W�r�0e: ǿ�zB� �e���n�re��Q�"TF�;\T_���\&��f��6���e�G���:;�i�����ai�²{��d�T,Q s5!sG`��c�VW�Ay|��}�,Ui�e�j0N��q�#$^BY�B	�\��.{��i�󉁵�q�����*�&)Н���&�>��?(kgq�-����`�:G��j�b�+A�ͳ� |�%�ńݤu���T���֯ܜd%G�t�9�����r�TZ8�� }�-N�]���?���P8�
2 ���!�N�Y��+_xĦ �])P�/\��&c�<�~���&�W����6����o�&"mlt��n�ϙ��mL�;X�8G-�T'�_�f���!g��!�
���更L�4�ܟ�{@��$fE�g�O��Z�M�[�d5�4Y��|�������|���t>�S���0�J!S�$n��6���66 �B�ax�Z�ŝ�fߣbc��za�v�ةA�q^���*�f��C���lu&�$��ݻw���t.<�>QEx��Ǳm{����4}�&syD�S�`��Sa�s�^��$G��J!wVU�*$र����F����{T�V)}����h^U��@�	@Q��BbS�b>}�L�@W%���8��'��o�C�I@c��A��W]�����S}��Ul9�d?0��H����-�
x���yr'>��uI���e7��b��d���uw�
��2R�PF!���-���^+?����ׅ�V�Ep�9@�l�=B�zlt�՞���#�ѣ�����N
�k�G,�I&�lBgf� ��`�X�S%O����
�����Tj��A �v�~���D�P2JطF�m�Ц���)eƣ�<���:)�z��D�l�K�T��%��n���[],�&��4=�����$���YLCKU�����Z���>CbϺ�,5.\�d��뜦�1��;p� 0,�˓B����2 ��	����յV ��)��5��4��5�a�\B���Lc:]7Go�V��0�3o�%��{�6�w�}�r��noDh�f����W'x�G:2�8)j���<�f��܎I�Z�s�{}������
Q����O�f�-��ȥdl��}�|�@�/�|��t����0���Ó�H��܋�
���fް�K�����|�})�V��ś��C~RG��jd��Ҳ�3�)-�jx]�����$��lST����'�}3����	��+��Ԅ#I��~@.KU. j��[��=1$��15&L�eg�����Ƽ x`Q��1�8P�θ�Ը�x���2�I��@u|��և9�(xv��� �\U�/���6�fu
��f㤥�am�.��6��l�����;6"��Ҭ��4W�{�X�M������!S�����{���M��z�&j�X� �-O1_�txwK�ٗ"���� &�,V_OQ~��oh�;�m��ߖ,(�T˞�.h��Vr�Z�j?�G�'���c�����o�.��v�,uc�$P���*�	_��o}�1������޼��:�)�:Z�q�6o��?:kf��L��5���l�[�l��fgZ�XY"WʵM��p@���F��@��.i�lS��Td-�!�h���62�>`EPN�`s3�y.L��фܾ�Unʥ�o��wHJ�U�`�+58_zI�{�n<tМC�tj�~/�m�X��]�Rs�F^-�Fn��HYc��;$�-�6^o�bq!�i2 ���GҦ컇�K���S�Z�*�h1?�M�Z�����y�KiG��RrAׅ4,͐�X�n"���ٻ�k�DUdB�I��Z�4�C�Kۿ�1T�x�/�=��˄����AA��:�������XU��owq��ğ�"z͝������Nl� �� �v�6G�K�d��h�hns<�nF�l,���������,���Sw�k@�sf�ܯ�D2�y�ͅ��a�(6�6��5NL�5#��:��=���=��G�����:��	�ܺ��c�kwx�;�m�SA�q���Ҳ�21�hp�\e���NzI�Ӎ�Oh��� CY��p���<X}�]#���mrҹu�$8z48U��3�#�:3�l�K�>M��{5:ʟ��_��r����U��I��k&�we4a'eٽ�~��g����(�t]~��{�!_j��X����v%�i�M_��ռ!" �v,/�dQ�֎��Z�P�'�PoV��P�T)�2�y1xf�O��+~��H�E٭do5���ͬ]�Y<�j��E��M��앰������@�_uv�?��]!��=�Gu[�?G�<�g~GfL�6W����ql�ym��tZh/7�U� XF%���C4C�
>v�lE�����b�+�-�"�.���@���Y��Arb��p��ߟ���[��cR���pQ��
�u�
�2��0�]����U	�χI�q/��إ�Q��*SWzg��E�D[D�m���Ɏ��pk�Fߎ�b�Al�߿�V6�H�o<���*�wt��NNL�Ms<52`�3kH�U�����U�mosn'��AS��ҏF	��٤���=�a���b�w�R��a#��#��֗(�k�U	�"ߌ�+����1ת���/�J�ӆ
� (�{9E�d��<�G]�ߝ�j�����Iuۯ=�c�l2B�̐�c�e����|v�isǟ���ו�o!�%ָ��l�b���4��0�|f��� �!��U>���w�E Y�}ǥ�oZ����G{�{�NF�[N8���Hg]�)����3�6B��~ԥK��Z��)�u��Cw���ǡ U,�Ț�vS�=���J���I���y13gr���0'^ V��$�Knl�T,z��$�}�N�w)���Z�7����� �ln������_��#r��gD����#��z��X[y�{�SO��S���J�X�`jD׌�� �Շw�H�ݨ���ϧ|�g�qu��h���
�C��5����wX�c��1��V�?��r׊9S�K&iG씉����)F  �\ۂ
��
�O�i���>곓(��j�-Nܥ��c�l����T�m�����5o^�z��ï�݊��KC;J�_{v�bl1��WsARl�N���}�^����Kp��J|�>�!_7Ș�Vmۯ������x����>:��ur�)�h�^�`���N����+��eS1W�1I�@H�W��	\^w�'�A��]��Ӈ)���\_�d����n�r�Y<�"���d�q=�$�]R@��O��N�3Y
9��3�Q��ɚ�@���K��f��w,���������}b��z��G�j��F����Q����4ݦ��^B#8��K���x?��%5��)]�X�ͷ�VۗjX|�S�1_�/�'b�`l�P'^�����<Z��}Cql8�c�����3��l�qX����C�F�,�1\ڎ�
T�Zv���o����j#a?�)�? Q%q���o���T���k�e���-$j���j�a¼'�~�r7�7˺>�[CQ�Nx&r��E[CĂm��ZE��k�>A�6 �a\1?��O��@Q�f_E��~Râ�����3�=�×�"s�>����I�YI�#�L��$�A:jZ	�Sq�GF��v 8����,K�)<N/Q�2O{�K��)�.#�����D�ZѼA���1:��_W�gV-ڪeu�����<�ʹ�i�+	}��<aֻ����"RZ��/�+9]"<��	�2H.��S�/.��r����A�2@u��9�����~�{�̟���$o�q�c��F�D�Ao��z�����[F���"�)j��C�h���yQY+ɧP*�������"Mw6��B�IcpGbJp5
0�9K�mx��i@����J���i��-���������Ύ���U.����Pl��������i�lq��>�>&�fG�Z]&�F�Z��>E��mu�����u+>n�3�*��}^�8���7b�X���N"Ԣ��:<����7f|�0���5���	�v�s��������OS˿�o��+��}�M�g�y�B�3��8�\@/�q�p�ڡi��me���_(��1q��$p��9��Q�+P�[��D�V�;��n��������D�3m��ɭ����[�k�bFܺ!/�?�?� ���~�$�����\�Tw�Q�t��QsȆ?�o&�-�첶�AT?��qKX	'��q+h��j[l��{��90���Ѣ-�4�sQ�Q�k{ ?�DEIS��~��FDk�,?#n^'AH���m��z:V��H���ߚ|��[}���t�ęI��	�!����������?���|�sh;�\��?ܤ�$���]B$*����x��$�CT����Ȗ��:�������?�o������*�U0�[2�:$.�}��U#���є�b#�-��)���j�1�|#�W$)5{��I�����S�3�!�Umm����	X�S�ԅ�^2c���p���M���>K6d�8�������y2����7y��p��-�ѐo�M	I3��v��c'[�@��'{ 0=9y/�!��.������Q����ah#�ʓ����Ң9��rw^&��޻{c�)숴�a����R����edh�f{�w�ޕ��eu�`��:�`�a�U9
~�훀�fP;�G�J����SgL�\W ���Z��-�L�H�fE�Y�CeL���P�Q���U :��_j���#�����RqB��惪n�[.� �v��Gj��<n��Q�0ܼAX~�Sdi:�Y
z*5����ޒ���ʩ��-�K��0ޖw�i&o���~��! ���1(cP���"J���n߯qI\�;y@�:q&n�mQ�YI6�Z���UO-�n�/,��B���U:'�]l4����\";�w䒤h#4�5=��L�!$33J�T�]iE��������D�=Z��ҙ��S�^�*R�1s�Q����P�P�1���gQֳs��K�* F���{`E֯tv�}����D3�� 
@o�� &֨-�L@=F.��чy�I|k�J	d�X�w)�0p�t�oe���'�U(�`��q�Y���_���u�;�</=et%!J�z���\!�x�3�d�%V\�*���#�f�^�"��SV�Vp<8bW>\#E���2z����N�@t��BB9U�K��97��ލ���)�<���WSQ�f!�D����I�`���A�a�Ȱ�g�N�p�q���1J�Ls�XCٴG;$̧X����� ���#/^��C���ڻ��٩��Ě����Pã�.vy�Vi0V��W�-�_��]�����,)o���2V���ꌀ��"�#��w�6�2rd{~@5��PPq۟,VU��l|�t����_|$�] Q�#�"e�iN�Sd�hᮑ���ј��mr�F�����}��!��`^��:�������?q�����Ŕ����lX�]�'�|r�M=��`U����{�}- �d1��z-V�+����jb.���4�(�b{��O�i�͓Ͷӑ�����5��G�;nų�XqI�`��.�d�!��"f7̃��a�T��ܾ�^K_v�����FU CxO�k?%B�ǻ�O���v`������!�fj�A�FY��(���.�}�|��u��Bx
S�yC�*d������y�y���������}5e� ˬrEG�LOt3]������Kf0�S����U�WI��<�����+�4�%�{�^Ԟ�8ʠb�����;�N
������=�Q��p�f����'��D@y7+蔍f~g��=�1Ml乌obأ'qN)����`��=����!���X�-+��@�O�n)X��d�T�ޯ�9(�=�;���4���F,��q^�0��^�x�;� �lH���'>���o�Z�p���*����}E�]]	�F���7��X���L#�Hq�L���i 0�(��wM���o���l;ɣ8i�a�?�av�6���oev<�X���Ųw�F����<�g���&�'����N�4�Q@Dy֜/�g�T����*T������8+(��1I��	ai48n������Lհ
|�@ꤨCOL���F���fzD�z5�ky�{vI7�0d+#^c�[�-������Y����9�5��OY~����x�rq��)W���b�e"�������+��'�G�͒e~�� ��C��T�}9�I.=�I8�9���C0���r5C�zϽ�~!>i�5��LB8�>)�{\��+�=6�z�<��պ ������"���Q���-��4���c�z�0ibX��,�����a�R�ƈ�U���8M���?��w�y6�]0�n_s��f��κ��6��p�V�R�&�x���Y� mwg��S
%S[A���_{l�����j)VUN�Nz����B�y�RS���6�}���V#�u���+��؉~�Ε�
1H�@�(�����<iB�z��x��Ǜ�e<6��X�� ��{�A�(�E:�`�#� S�&�`��,���BK ��-d��+,k�B		U*���	Ս2=H��f�
Q�q0Q�1)ռ,�yU���U����͘5��tcM=Vqպ��;Р��%���d������w��>�@�:j��vQ�7�0J�����+��R�'-�ť�Fu�8�f����úK�S����E��Al5�d������W�l���VǲQ7�E�b\As_�0!\ة9��, M�㟦�^��z�w�	�dYY���wR����Bł[��E��'�5�vR�	����m=�Hᓫ�s�e��S0>��c4�Kh��ok�E6X:���㹹��bMi����4�� ��`YE��E�~�i�*�$�g&��YU��8��.�V��[����+Cމ��¸�T�S���ܱ��{#�≸����тJ�P�v�l�	� b�{g�� h�{P��RKK?�U0/��~��W�"���FH�(�*�3K�$�?��׷��`������7&g%׻����S?�ؓӡE�[v�[Fi(�	l�zX��;��8��K����A_N��Ϲ���[��q =�7�vt�C�U(E-�	#��ѽ�&>���dޖ�V-�(�)Ar��)D�G�WfzP�O�U׀Ǳ�����X��H��KQڬ�+Ԅ"v�P!�#m��ó�pb҆��a��J汝�/����a�j']�XY��6h�r̚�pT߬y_�LCpA/�F�rCE�zB�h-Z�D�Z�+$�6�f!u�*�l]�4��!M����py�!�$kL�3���z0
�L�Cn��W�ޖ֏�՟7����ku�p-X>��`.�Iª[[��I�ă�7\Q%��c��ޜƆNvC�y_e��N����[�(�9he���hk��#�0e�1ڝ�i�c;,��O�W����}ѭ�DHvc�Fܢ���zs̚�:V�^�P����X������m���R���SO�H�GR��	$ԝA��M�廆e;�^+�,6XǓ����b*�f�o���?a���l�t��(��� f�H��>*����
����^�V����rP�����" �.NF���y�ｽ�������]�J]J(VQ=%^�ƕ-�8�?�lO8�7��˸.�h�=<3�2���7�O9>.�����mF|��*���9�uY��ʜ��q�9|�X�:6P�k�|Ʈ�d�?��;��ב��^�c����7� ��aGsU���j�4�u���E� RYrW$.,�'�����n3ZTzj������$���ڋ���{����f���W���Uw�FM�ÈJ���5��|fK��-M ZWn*�K���'��lԘ�r���_s��b�1`��Rjt�^(!�d�\��#Ѝk�s�
r�)�E*�p(�}�z���7U^�,1�lQ�xo(&"��@w���1�:�"��̯�H�/E��/܂ Z+a۾Ƌ�iI�˗�+o���T|׋CmM�K;+#5O��jɆ̤#wy�Q`��A�<� ��P��Q�e$��_�ۡ�t�XȘ��� -�t��'����\
e��&�PU��ɿܦv��e9t&tX���I#' �:���Ó��a�j����4d�_Gu�v\�`o���;녗]�D�\�OcU�:#�D�0���Σ�> ���r�@T�h�x���T�~���H��:u.�6l��7�o1��Z�Q�H��V��J� X"rr�|��RS��=wq.����dtܐʃ[�3���{�6�@[߳�sj�	HD~S���W��޷+_�!��t!))紿��Qj��1�~̩�U�~m�*L�H���!8w�I���W�����a�CX;\#-�Y�CSǆ�\�� �20b�{��j�f�;;��S��A6��Ы c \���]�ƆI*s@ U��{gJ���lsߐ_�}��1��K20��m�#մ���K��s��\)
p�W����ъ�>K�(9w���F ��d]Y�>y��������?���{X3�Q3r�|�^���y6������Cg�q���?5��Ԗz��*U�\	p�n�o��$�38��y	��.R�L���j��1i'8�e�<f�P����9�.�*9�2[�N��V� �8�z,��kʾs�|D���U��w�"5�v0����q��{���i_޽��.��v�Ij'�uY�63����HK��҃G���p�k�1�/e/��@�A��xrV�k	,�r�)f�3�hґU��5H:���̱��� *�w;dz?�	��20���-���޷	zT?����s턪��"�˲t��R�k�>�_��-��o�����/ƻ4�$N�X�=�r��s���b�-���.�!�٧&Bw�%{ť2�y�R&�w��g�o��.�hx�ڽص@4g�`F]�B�0���W�{$��X�S\�9~��9����A4ӹ�~���qю��0�q���uWĎ�+n�bl�&�o�p
���z�I8g�u�?m�֤4��˶�r�=�������v��L.'[B�k�{�W�����m<�����je�u�2Q���O)��[ojj����z���'�_�<Ȱ~`����-�l������%��y�&�����޴���N�-I�y4��ty�Am�oSS%r�s�$��������^�>9�����#X$�%%l\vx�0�8�����[$���[�����A���$�b4Ȩ3��^���^G��w$���dv�����Ï;������B�o�l;�d�>�;:�\-��=<v�x[zRX�`׽қ��SУ�c�e���`�g����UQi��n+Ka��Fs�D��,et�U:��-�y8��w�H�?&����3��I��f��ȫ�9���?�yH,�S��Q�����¼}6U�2�F6Qi�v<�����ݣU���O�AOJC$���,�ԭ���Ւ��Aj��?/|jl�������6���ױ�`#�&�8��F���ٍ�T&��k�i�V�M�G����4��`^�9�JݧrGpQF��@��:���un<;<�L�=C��j_�ƕOc��8�_���z�~)
E��=�awQ͞�e=T�1�ktm�i^�²�2'�3��3#<�G�^5�/f�k�{�.D};��!Dvf���^��n�PSA�(��}�XT��-sh��sS##�WP��g�ĝ:�uP���� �T7XW���{�.R��m�_f��^�H�_3�����P�k�m��g5=t_� JEE�a=Q�1��j䣇V�)��gݱVx�	�W��k-�{��C&ē��͠΂�+o���C��瞏����f3,��r ���²�3�!�o���i��d�l2��,���ύ�E�2�5^D�P�Dgkm��E��Jsw>~�
)����]��s��Z���Yd}y�5��D�y �3JC��U�����dg;Hһ��O���w�W\�`��)'�˱�8�ʾ/���ל�?*���ힽ�d��R��M7ڀ��� ���Z�7�БI�q�rh&ScX��GyQwH_߲���2Z⌣<G3��@r.q�"%^ΒRς/w���0 G�7k$�MK��:F���i��֚=%��]j3J
����`�c�gW/�T��FGK����2�sSz/��h�h�#�+u����&��R䷺�ioQ,�\�?�����^r����aLl�FjG�2�
�-�S����:��4��Q-���HX��#ct�k'�*�$�dt{ =������i���e�-���Τυܟ
6���Y�EI�|<�7H�s�^^=�����Y{�Q���٥����hVFv9�^u����C<���+�3mڼ- �������9�P�S��OTі.W�0����#��>��Q�����q�S�m��5ٽ_���ߺ�5S"��YyP_R�jZW�/t@��s�F��0��k�0����2
��� 6�L�O��c�҆dH��E�7��h����>���-^�V��SLd�r��������Z��D��7#A����u�y��^��}H0�ҦX����<����ڽ/"F�G+~37 �'e�9�A��`8#�_�}�Ww�X�����v���5��kd�%�AQ�*.��p�A�6(��������[�N;�W �!3�h�(���s�~��<�i�%�[�~��R�_�O��)��*b��q�����fY�_��&�.��t������Q�REo�`I��HQ�a՝h��N��MyꃺK@�H���X�o����|��n�bD�8���m�zl"���6UkVR�[0�'�'��ĩ� /�����c��YsĻ]Bx"����WB��]�� nw��9��?�Х
����8n�U�F�A0v��6(��x��*��#���}�3����p�n`��=�A {�-�
F�R��<�YP�ɰ������ً,�8xw�e�W���X_���V�GX�)���BnXt��rl������vf�JZd���+��"���r>���� �%�ju��G�:��
A�c|v�_]�(�K cԺ�	���V��B!��ᙇ�����9�,a��^,[�vjޞ��`��h� &��iq/�Su�}&��<����i䂹��}@��'�.ט�fm٠>F�m����N�V$�x{}Y�;Ɲ�|dc�-�]�b9(b"Fsq�1�
���-�F�_4��!�w��g�G�V�.��$N'��ζ/��U��%�v�iK�4��y5�u���TƔ���	��nU*s#;M�}�5o���F��;�NE��_t�C��s�b�{q�*���},d���+6��L�^����U����7+/�*�{�K^X�E��?۠7�� ���pgp�i�c��oMMF���"���5ŕD�O��A��$������W�Y2|P�x���ÙG	�G�h��l�wV� s%:<)~u7/~�}{��A.]��G1Y��Xƞ�P�������G^8��m:<�3U;���җ���I�>�ny{scy��|�1��7A����R����~�����̄�,�w�����[~X�[Mr;?f2%=n���ۏ��Em'�p8�V��@�w|/#V��3+d�8u�{ڀ�t��Y�?�`T�9����_�[�̬=����\N\�Rip!�X��*�V����]G��Ta]��[����e���=�A���7��ŎotK�=���z
�h����h��޲�a\����TB�����cq��0�_�-3l7@!�u_��K+`	sO�x���b��l��j��b_�K���75��V2����	e
jd}"���-O/ZZ�?T�ڏ�XqR
�v,��0�0�?���a��t��U�����5��Pa��d�p�[�66cH`nU�E�#�o�هk��jt���;V�"��4�D(Ollchwx83�<ަ�;is�r^i��xo���:F�����W���Uy�S4��Z��/ؕ����,E�;1������$��]�2WLF;��b"G�3�}�R	���>e}s���BٽU��Z�ԝ����`���c��nz�c�:���&X%�́nɨ�]0���P��r�~Ws�������r�"�@H��,����ؑ�$����ц[���v|�4��*-M��5"հ׉��e3����g*?��<��~R}
;�*W�z̖!d�=Q�C�c��x~��$ǡ�2��:�T���8��>ILGI�@ ��Ը�kz	2C_�"�sǰo����H]zN����/#�@VE����Eќ���K"�߱�/�~d�u �]�r0�7����i�=�<	 ׶����xC=w���H�t���>9�[�5 �2X8Q��^�E����,���!���$3ɴ�&������o��k� +������
2�cZ[��*�A��b_A;�	>�q�{�}�z�݅@��〮��mC I"v��Q!>4�ˢ��b�]ݍQx�%3��HB�KƬvG�^Pd�_�t�����؅Cx�\�$�g�9{[�]=|�2|k�D>���5�T�(��^��6d�щ!�{��h=Vyjb���N*x?Ex�^s�Z���e����ֵ5/*#�46��;"ʦ\\�6�������X!Y��쿛���{qD��z�)̺DT�9�iʀ)�*=6��@۟]�x����i�>�����*��NЭ�H�<L��H��xKMm��&�#h,�F8��P	B�A��0��(�tR5���(���X9�$�Ĕ��kl9�<sW�*��k({�a�W@9�K���Ϟ��3~yt�{&��2A
�ۗ��U��X��Ђ��lT�!X��[,�7��l�:�� '8cb�v�K�c�sBLF��t�y�ZĴ+���B;�O�1�ˡ݃޺�o(����蜪s�2�.o��37�ҍ�f���M�%�0 w�k~�F�9wq&m��&?�+�I�QJ�`���ޡ����ӆ3\���/hX�5���>��	�'/�"'�D"Jm�:�SvB�s*�
�Ma_�ƛs�u��v�R���p�c3��;�%#����L�"IKR�ō�+gSkG�V�������������qP�g��q�pɸ�|Ȓ喁�S��!Cn��g�Qe�k4���"O�*�q������7�Q�9b��L�8<�D��2ٵ�<w�F�X�W0�iu�lXO{J�QJ����$�.V���@>C�G���$�gޥ�{f\���ן�'���@e����K��.j�@�L��j�!��~+t�zǆ� oA�ǹ8':�b��N�V]I���J9�LA��tq��MH;��ٹ�Q#�˔�<PF0�� L�h����h�ۭQ�.����1�K��T޽|]�d/�w\A<�uE��YD@����[���Ƕ�g|<�g��TL�<�-ȿ�\�
�(���%+ٗ�s�+��8Ot��h|;�DqƔOr�B�@�����9F�;�~�UdU)�2PBRl�TH � �3��	�k��"4�1:$�/����Ҕc�ǹ�B7�v������*Љ7�� �e�3y!��w!e�H]~r��0��
Da���A���T[�h��tg7)��A�,�X}v���3�f��݅1J  g}�E.�#q�5��@K���e߅�@�å�f��1����u!�7|��<Sd�)�p�8���������p�[��[�����rJk���c�"�~��O���OrIBp�m4�s��j����+��\@p��qiʸ�����h��]�.,�N�w
�.e%:f�!�a�VO6�,�RKN<4O\?Nǃ��ȩ�-�$�|(ů���������"�����V�?�(�Š�q�1xXE��y��L�^���	�L����d��;)y�K�V��(��If���F��ZT�^�'���4��(�r=����L��u0$��9��>�_D�v�WE*R$�9��������2�ϕ3t���͉��&��x����nU���Y�u�dJzS����ޕ�~q?��60N�� R���U��-�3@�f�a���O�WrHI��K�#C��G�W$�f��~�}�0b�/�P�L�� +�kDf��<n�4�a�	�*i�H?44�ݭ�nK���U�ˎ�[�f]5�$�������K��FP���/���A�s��[ |爄��e� v�B7)�XYiDy�7X={��IV��j^ğ1�=��?V-[q��+�����w)E������nȓO�h4F��n�@� >~��H[���<A��Қ$�	��:�𙮶zR�xu�ɽ�}�<� �����1E0��$�T75��.�o�]�A}	è�#�g5ߕa��Z��x�z"a�έ��ZR�YY�tj&�{G/oe��@8����"��ሒQZHQ�
^�Fa���~Ik���8�%ʶRA>��!qT/\9�6^���V�8q��#\�vX����B��"��Mo��VPx�U����;�s�g��r�^b���z��^�6ɓ�c;}���eԫ:ʻ���O"P]�b��D�%k���U�b�.z9J
8�R� ,<-���JW��6F�
c@o��o��m�X�U:s0�HQ��E(��Kz�"zdiI ��#�R>�p��q��A۴���6����t8Y����Ćt�����ԇo�i����0:���[���ٔ��b��߅a�	�9{��@�=���d!�h0�j�Ç@�2�gc[��O���(
��Pb�?կ���O<���;��cj������= �%g}�F��א�C�ɯ	�h��~t���t��w�j��$�eD9��M�R�G8��_o�mr 0$7����m	i����N�C}��y�`� _�K��1E׿�3��RHG�Hx:Qw�)�"��)�^�{���gF����4�,��i��� +���S�	Yc�C�8�7�{*�:B�h�I>l�Ja�~�ڎ��Q&��P�,�-��콅������C�ry����`W��؏�Sq�������]���O����(��k�و.ǺfA��Ik[����~v�fX�� m|ہ-'qϭH��?�ZcB�d������T�Ѫ�����ˈ}�x�\(�����n�r����tm�G2G�&d��A#_�����l�՗�&CL���Vy����H��>��J��
U`h�x�_ T���M�%�A��*����+[|7������Q����G����w4#�n�C���&╮8��Z�Qas�k��*2Z,�`g��(%�_P�^%Ŏ#z��B˂�Fsو�Fe�Zc����T!�^�d��(�u�(�uV��5f[D6Uj��,��v�]9�%��25hn�����X��ȈzV�i|�$8,�Z������.�k��nj�dL�Y��q�6=���c�\5�������[`û�x����*_�Ԃ�yJ<K��	b�����B�\xU��F��W���?i->�%��)��bÕ�4��S�ʹ�s	���T�����̱y�� ߿Ͱ��<��(�����Ż� 4�8<R���:�蜧O�4��G�TV)-?�N��:]�WHz�����G��m��_�;rx���l�s�l �Eڊ��Q��cC��cԾ)��+��h��my
�t ���3C��ec1��f�`Ƚ���P�GK��'�G
���N��0[��Z�(2&|.I��Q�;��e(�G2�^��+�Z�el9)���.��#g$��-#�z9C�X �>D�Hȁ�XD�q�����7���7g͖0^
�)>�T҅s4o���%��`�^�sX�o����'~#��D�<|��U)����5S��uI��3�+]|J�A�ꫴŌ٠}�3��Æ��c���D�*�\�J�I%A��(�f�ڤ�,�}�/�O!�����Z�\\���싉x��Bl��1�����d�$�D����K10�$Q�LǟM��	��T�#f8�4��)�gs`�I8Y�*�K<�ѮJ������N�����%k��������a>F�}�K1xC�We���͒�%���)����n�Õj��:K�C�.X��T���`�~2�ʓ��Z}+�ܩԩ��l<�oxϓ�u�~�H���l����%���|C��c��{�}��k���l,'L�kE5���+���������^=�Qx��<�K;��G��/R9��fh�ӒG4<���̉`!X��@X�'�6(�D��˓�Bʔ��{&��㖉<�_��Yi��e]��>!EмV��˕�"O�S/��ȪgJ��q1��帀qc�m�_ïe�%���ʩ�G|I��n��$���e�ۋ�P�7�S��<Lɂ^�	�Ǻ�i���4��p�r�>�:�[)�>E݇�j_������W�h&ɬ�O��P>��ϝٱ�iEx@ƌ\�h��XS)w�*p���E�/��%%��u`��m�搧�|+OE�n#���"r��n=�ꋶq1#P�l�����O��Tn��bqI�V�>M�r ҷm{į�k!(g��t˗����H�Xm���`ƽ�����l�פLB�du�ȹ�|�D����o8|m��q��	N����8�b����-�E�$U8�����oJ����R ����:��/cw��,WS	�Ų��$�&�b˵���B�����ѓ��g���"�_eN �+;���Ό��a`��(CJ�1�n�&���9���O"�u�2��l!PJ. 5ٚ�?/{!��^��Ϥ9Jk<_ڣ{�^=jC:����S`Db�O���0(eu�RU���o^r<eB�8~�-���Y*�5�o����+d7|�Y�|_�_�|���W�b�/Ҽ� �`qڡ@R��H��"��^K
az�~G�0�����Lޜ�y��Q��y���(b6�bI?Q9_��9�R ���I��'qmL��V����
���At4�x �*��a�Q��|j|��*�z5�N�W���}Ъ�:j����46���s#v����[ӭ�os������f&���L,�qf�26�!� r�A(�B\\]fT?�Y�_}O �ěY��%Ǚ0�2�K��35����K|�RA����w7�t����v0"�(ǧ�,�#ӳ�b_w���ߺa����qL���jRH��R��,X]�q�?�6��}y� t�Օ\X}f�[�u���h�C�*��u���r6���f�gA�DJt��dD�����|A#�~�J7�L�V����ۘE�7����çD�7�O�܅9o�(��ɻ84�\W�߾�Dc��}Ϙ[�S1$Fz��}��O4,��-�Sm��M����X07��dQ}E�i�b�쇐b����sIYV�-ZOu&l/S��zCY3����$T���O�?���t&�l[A�DF#Ss�9�6�[�%~��V ���4�
����ǩ�OZ%g�*������~�Mq'��@�m�o��L�! ���/'�]�=<>#Z�[n��]�8��<[�,��k�	ֳg\![�OÈ@�MIN�_��Hb�PJ'c�P� �!:��MT�J�Z!�������.V��cF��Mm�u�O&
�!V�^��2�����^�Y�5=S�_�}'i7���\��Ҵt���]U��!O3J�@��ě�#���g��$�yFI��� !#J��,V�٣8SxY��!���4a8J}#u�s�9�3+&nXD�����oa�?�2��+y��*�Y�DХK��Ƈ������w�������T�����}��$���P��������E�_�j�Ʌ�>)%�H�M�g��~��`�v5Հjʍ�&�3bt
E#ݠ���M/���`�D ����2؟���c�!��P�ko-5�d�U��^PwSVP�������l�z�4�>]"v�4뼒�bd�[N&���eM1��7���T 'k�v��s��AR��|�|����o~R�z�;ܪ]�ZM�~�ا;��  K�װ��v���@�f4��-Ƽ�{�D�Ȥ���u{ "��Q�8�u�|n
��R.�B-� Uo1,��T��ND�~ݎ��3������@��(��=B������!a�����q�t�HM�S���iZ^%+:/g�=`����a���Eu1+;����<�[��`�3����g,�_h���6��;�<�6U��ou�e�Gg\�>;X�LzȈi�'P}Q V���d� Dr��*�n����۰�b<n˕��Q8�ţ`2��n$�W�Z#W��+E�����K�:{r����jx�sP�/��pP�E�9�Iwϻ������MKW4=['��䲛�'q|���v����0�M�V��6�
1�������w̴j��C;	���؄���v�dBx��<Yy���0��NA`�@�=��Ώ��s�l� 5�{��B*Y9/aC��L�o�ڝ]�caDE�1����K�Y�/�F&N@`Ȅ.�K+�󳬅��h�K�j�Ȯ���H,��C���%�pM֠�|���t���1M���Up~= �����/I��%O�>����LjN@���f����W���~��B�|�)~B��,��0|�3��+�$/B�S�Z���	.fC@�'{b���E�$��ne@@��v�������oH����a�U��j�ڝ����*Ua�'�ݰj�3f��`����q��	P��H,~G��
��q�y�$�J��e��̄A���/���<h�*PV��4�Li&���2��^��@H��u�%�E��!��<�w�|�J6�������YC[���N�t���X��P��n�
�N<�#@)W����������L�����'h��JvJ��P��~6.!n�)5��dt�2�=*�ٖ[j���k��]��Z��T��q)��o�[��+c_-D
������uo�cλ;'I�|�L�t��%���}��T�(�n�o7��6X���#?�Ka�RN��׎XB�nd�~;trjȻ��H����,���>�Ay��ED�ɣ��p��J�7
����i�E.1�Y9�I�	�-���T�;����	k.��ͻE�[��a㜂^��C#�T��f�R�̯k�&���y$�U屮aI�w`��AW�X�݂L�O��O�¦��&��t�1(�g(����m����Q/��Q}3��K�X-�L�Y!\�>aGb}T��oAf���WhM��(��ϱ� \�j����'lb���n��h��/x�\��z�%`[w�$��r?�%�/}�/5�$��B7V�1p��;�t�ず^}F�U�@���9O�'�'8�iR��p^��}av��Uns��e��!΁���B��:��f�[�+XV�2&���vU7���ލ:�Z���@���&)͋"S?�'�B^}�xKƑ��=� -֠�~�.޸'}��e#��	�Ɯ�ʤA�����Ѫz�ĳ<>���_�ޫ���b����X���-�׼Ѻh�B�6�����Y�M���Y��7�d�rD"0qn5Ot[�Uv�X�֗h�)����*�h	5/��D���;Җ��i����qƶܜ�"_�Cg_��O�U���J�T��_����1�pF��xW�`�0'f�VU��t
�<�9����о3u?Z=?���3Y����!�xb��h��:�R�қ-��mA���Ըl�(6z�}ārlC^�z�0A;O���Z�UTTJ�oe��'���BQ�P�N�jJ�5����u��xKY��z��q �E��9>^�P�K(��5�n�9��$���1��i�M�M.����0-�i�`�H�Ili�.�2B��CX�sF���^�-��/~{c���.gF��lX��X��&�� ���z��W)�p0X4��G���,3u�uD,<%�O��Iv�bL�����hGHz7�$Կ�(ict�0�n��c\ȅr�B6w)
���1?i�f����C�7{���c4��V���,��%^��~�������=�O�&�#�P����)G欴�h�X������:Z{	K�fdpPm�,B�mU����2�Z�ݡ��j��L��c�4��4k��GŘ	�rd����c^k�cLk5�������z��>����錺p/��؜ײ����x[�Hy5�%�uY<�^Fy���0�<%�4�۞K�0ʾɍWJ/o>l��� *�j�
T��	ZjD�ױ�.C"j���P�1���V5_�=MK�h��Ǹt`g�F�oq$j(�>��6%���	$��;yS�u� I4������p)�͆[���b4�?�$SO�FM����Ί��*(� 3:��]�UM��XR/[ڒ b�3M� �f�Z[*�����-d@|�L��m �T���f�ٝ9��?+ʦ�"}��N��g��u�k�i�48��q�<y�<J�x�������qL@c�K�>�疻�D�eat�yo����5>Ф�S	�T��z��C��K�y�������.��fC?�g/ʨ�Eogҥ��5�S4k�f���R�|!~��R����U�)o���G�G����	��0*��r�x��mYgm����h�e2�-�N8Ѻp=����r�;��̥�dI��_�sR�M�5��+-�,�/W�˛�Fn��J�@O^�bD �:P,m �Yg�=��Wz4����*�#O6�:
!찝#�.J�ր(n��劅ob_��Y��Y��E���iY
���H�>�P$E��ج):_7��+�����"���QfTz:��P��yO�oimw��6��R��Ga�J�7���s��57��>��@�`tuM�aGZ*�C�[nn7)�E�`��q�ע!�.qŏ�7.*�����QX�'�����R��t�/A�}�Ml��KS	l$�d�����~0+S�0>:t�m�7fd�!�qz��%�g�Ì�d���2XV���Ѕ^eh��orz�1��m[)��\�?�[h6���p����iI���S����p����J�{����u���o�lȫ�UP�k�5P߮u�X�����{e\�ʉ��<�~�p,��}f"��;J~eG�O��^����w5,�L-�,���¿`[�2Օ~ث!|�3�%V<�M�W���/�\'=dz:-~lS�3M__=�1�i����_�ɆF�Q*fW��:C�i�T��U
{��b��i�ͫV���Uu&�9�����I�PīZR�u�K����W(����1�������%�"��@NŝV�j
�0�i6�Q\����/T�m�N���%
�&��@��Q���#�G�n
�B@_.@�:0jt�*�ÀzN�w4�5(�m�]D�
t�y�b��F֍�x�aHA��,N�E��+����
�X�Ѱ�s4~@�����F�r�V#
,�� ��n�:=����8�~�Bp��'VY�\�VK��by��=�R��'��Ma)����+�����Y�C� .m[�Z�D�*���I�b����--��X����S����Iy�b�H%����@V��g��p�T�9�}M���� ������9�&R��!�Yći��w�Il�HNT�}o���@X�;��h�|�b�~��g�'��5$:-N���
i	È��	���id�h}cZ�2Ѭ�-���Ih5eSbR��>t@RR�MP��1*�';�4�[�և���QT�lx�M��j�JŮ���-�!�1�4��Mv�~Ǣ4���#����GK��Jn=N\��Pjʣ@^�m嫊3���6=�)�T��V2�%�:����+n��'Z������Oz����f}�n�h���22Q����[W�� c���h�>n.[J`�V�{쀚o�����ѐ��XJ������u���oz��yV5��#0���7g^n~/�"��g�<��C�X8��c@ V���T�%���@~��-�Yʂ��ZW�����K�GU��jsR��)���Ԥc��7���o�a�s �2�ն�`�OY��`�T�;�W�U^��'PR�3ͳ�3-$���� �n��;�̕Īx�!E_r��*���n��	�f��b�'	7v98��o�MQ�����)4*��QY�=�l�(M�Z-��q���d-]߄B�
����J#�5���寨1y�o�7q�H��:���Aٖg�@X��xbۖ/A.�h�R��`@�5�k6�E���]��G|N�5B�H��|��5d#;����^��k�^�A��!p��M�EXT��s�pc�A\���M�+}&��ΨF��lq���9�R�5��Z�~}�m1e�}�|��?����g(T�˔^��e��ӂ5n�aZ2)��%*��]�ۜK�n\G�������u�5O�^�}�|�,S,�|�5�qY�c��M�SYo�l�9��os��&�7'V�Ǽ����'vw���7��;�+�=3P�/�u���t�����AL�0�e7�B���nM:\�j<��^�3a W�5kE�(��RGz�W�ջ�`��۴!��|�L:|eل- �n�k��r6n[AY5͡�a�{�l�
��C
��"
E�{���Z�2����QZ�^�"<(�
��f�P��O��l�K!�x�!�'�B�˓�)Oi�8����瑟�b��oWS����W���_*8?V��F}�d~l�<K�f8�����^?��l8e���習/F��홠�J�s�ݴv�x���J����֟�S��s�Z	�×�9�El/��Uf�|�ň��(e3a����0�&�� [C'>���am�����$S����%���@�����^ʝyַj/�P�� �I��^���uN��ӌ�;e�f���{v��eϷ�"N��f����k���)�x"����1Da�GD�	T��X��C��<�Lļ ���	���#Dw�H�\QI��k�T��I��]��
�]1c��Y����u(5X. o�Ĥ#�s
�$D�^FrD�,��� ��)_�I�ܣ�P�{H2�|/%��	�W�t�S�<���q�{��71��᾽� W9��萶GÆ���
k�BE��|h-"8�d3Hg\Q]Y3�����Z��e�+�O�erW�ޔ!,�����nV9%}�baT��&X�{ZI�>���_͉�I���u���������B̽ ��D��EH�P�c���2���GF�6��&���#f�������|�?R��ov�wg�DJ���ku������ɨ0s�/ �� ��9h��|�t���<����\�����M�������x��1?�^F��?���Ύ�;�a}�F�胅�*Ȝl���X���%8~��5�q�b��s���4+8U�X�>� 
yh�I���=���IA}��P��х�m^��� �v��^�4�ް��?[�����C��`��5�x �\�i����-����FM��.�L��*���&��Z�LD��8Y����K��\��:�
Mp0E��
���t���p�{�}L:�g"CF����������-VW&o���U�Ǐ�ۍk��O�N�V�co�l+�y���_j��V$�rR}\�!<�������R`�D�����)p-4T����G�'�B�En �����R��1�X
��p'�0-������c��=ohHI?��N��Rjl����0Ԑ� 6@�;� ���2�������������T`c2��$�˼ʿ.��.tT�C΂;q��i�|Nۖ�;Z����j���qE
��Dʏ��DU)��Z���ʇ<�e�6i[��oH�u��c�Oс97)�vW5t1��d̶U�vt�N�ja)�5���	^�C����@�Pe�+%G����_E���Sm�sr��*��UCT�М�N\�$��&��k��  ׷�/�n=W\WO�� "_
c(@�Ĵ������C6��ү����s8�pÿ�D���-��o���#]$g�պ	��@-d��QclS�1�)*��zaw��cɲ�I!w9S�I����)5揧@��
A}��aKc���N[��e
�1�H��"�C�Lw8�ӿ����uB���<��h;�����$ �E]�>��6��I?�s�Ǩ�F��\rR�����ۇ��'�ֹK��u1+����?��h���_���KGʇ�g}2L�Rd��i�]�#�2)�
���q�}�\�hS����(�.�v�u�0C2RE���%��@�l�$���S���#� ZT_y�E�Rb27hW�ti��H�������?�������s.��Z��FV|]�\�G�ѝ25w(-\$cC1�mV�x�N�E��ܿ��T��W���׾ڎ�q�IU�[�e�}9��A6=��
��+������T�#��
�~����z�m�����]��]���(ī�h�(��@���@�A{r���a�}O3(c�>!���r�?��a�X�c��rz��lR[�E�B�ZmV�H���ɛӮ�F(���
��%�Т㋣t���C�O�V(LG6t����Z�:���Iw[�8+�W#���sy����y4o1����H#w�웶<����\�ћyT6�N/tk�b���)Gq�yv�����:|��ԙ����ɂ��b5��ޟ/ {���'�Յ�BT��g��k�۳�HrXFV0���~}��U�Klm�����iG)�e9�Ђm���°�u"  Y��j��m�;[����Q�����Q�
ޙj"�&��1��,RH�`#n�aV"��/6��IW���57�zi�w7`o�o'���R���,���U��-���=/����y4iX����.~B�,�D�<�e!#�s��S���r����0�ג:ݦT}]CZ!C�Ӳ�[�`�=���sY����ih�zG^�z�4���u�T��je�D:�5�ݭ%�O�mǮp�v���2U�Dzx���\xšFͥ�ӑ�/��P�n^���x̸%ɀ��+��a�N��~�P�v&4��|o��̴b�2��oXjJ(5`�_��ٳ-m�*B��%P�?����!=���G!\�*ΖE:{��Ն�"�\� .R��	O�wz�L�Fa���h�Q��t8���p����wEw�-�5��kۡ��	�0����-�DixEn�k*@�:#M�9��0q��l9� ���oO�\�����/�7��s_^�Do�2e9BjOt���'a���B��n5�h%�9&�`��&�t>�:U���OL�ʣ�
�p�=�>�}��@f|�M�pC��"��'��,^R�8�uU"�{Se�j��(��25���V���Z����B�����H�l≺FD-(��q����9��O�O�V�-�%GrB#{�r������l����exO���A�;я�4��?z'�`�)� ����!����}Gd/��_��ҸG�w4�ϼ҃P��y��XL�&�׌1 fctK?#x���,�Y5b�5X���e&p����s��Ǣ˩w�<(^�b��iW�/lE��=�o4l�lz���ԛ��8-��M����ϋ8E�&�vP�o���<^��z���+",��-�V�@�ǹ��%��E�S:����A���iwk����Z� �+�n��bz��B�E4��'{*����zf��Ҩ����M����?,˪ٮ�`�HD��LZF�$�9�ҳX)�qc���S=j/E�ɟv2�HCihMb�4�6��Q�&�9���7�N��]1k�4���Sp�V䇸t�[�6��zy���؊�����-w���**�U���):�	w�]|B�J�ω�}89�)sD�!�^\n��'a#\z�������s��[#���� �B���k9�h��7yh����e�ҬFlL��9��d+]9ȫ�ft#��FY�4��ARZ�¡ň����Q���p�e%V���)]� nx[[t�o�����=����'7��>��u�/����;1����x1&C\��zJ}=gs�܎�U�f���;�4��k���m���ۆ��"�@���C��+�Ù�H� _��<��l*˃�T�5����ҏ�t*xX�LE�������I�d��'��cU쵍1�~��E�5��ް��Oܣ��*��`7"��ϴ��/9�e������-������'��� ]VMY&�]T��'�Sȫ��}��tL�*[��&���ly|A�@Gȭ������v-	l%&XMe6�����7�n�c�3�NSh�t݂iv f��Ժ%����?#7W^*,���V�_���l����ʈ�h=%��NQ�[�Zly����* s��3�?�8�c�Q����S(��EwE�F����VL"�#���HX� l��x`8�q��-���G��^�׏�:1��ezw�6xm�K�)�`u?F���w�K���	�r�a��os��'�:̍B�C�S� ʫT��h��q@XN2�`j��$M[0���	޼��C�tߞ��ƘI��̍
��n�*ˎ��M���҂I4�,i��p���������&����;�;�L���b�H���Y�{W�d�Z3�i-`��I����C/�����z]�A��u�o�^C5t��A����0���������X�2z<��K*�V���av��v5%+�@��\J�uM��/6}Q��">cjAP���Ś\Od!�m3�6���ok���o��+j���ٴ�ۖ����2]��$*k��6é�����>)����c ������9g�Y�Yv�k��-�5�0-�Kbi�9��Ư0�c�܉h�� ��qٟ6�����U�`�{y
FZ�qs�B��@����*�fY����xp�ﳯP�S/b.N��Gtq�+)�v�A�&K��Tz�!~�fs�"�_2dP�Se�+kg�����N'ϭ��ε?å�Ē������P�"�՘C�p�}���ӫ����.�)C�C����B,V���e�0˨ڹ1��^������ƛ�R'��p�X��Z�n�\���(��� A��c�'��8�isp�C-���F�f\T��j���)�p�g#���S��۞�ĖXj��k)g$���5���:�:Wbe,��h�
��ud��� ��B�kuj�̤;��w I�k��gs>WʤL[�|�8�F�>v����>��$@�3�lP�Tz+EAڤ+�d��/�H�
�f� �Z<�nq�spK��s����������pvȁ�fV��3�4$a0��j0a��QdǕ#����+[��Pk�aY�<���R�˓k����CKʺ����pv�����'m��U��H�3)���n��Mrm`4�#������{�(m<���'QU�2�@�(|��*���������~�3��<�it�-:�=�\�Bݶ�V5"2�����'�����}��c�3�(kѲ�-��_۵*[6����GX{_2��'��? ��Vh4�cgF��F���e��+#���7Z�.����pKH�3���D!2\[�F�z�U�vʹ��⶞A�Q4UZ�Hޠ��s��|Y$�z�5����X��W�|�$��뽹������03�_w�^u�G���ڐц/���6A��e;��Wd�%PB�~������	����b��rv#�Hf��Y͐��B�ڎ!8�,�f6mv%O��g�,��nhr��u�1}�Ӈⱽ��$U�[�S#h�Bܻ�}��?n�D�x��,K��Q��m�	��7���A50��zf���]ˣ{UE�X�K���ҹ>N�s@N�W�+.�V��n�"�.��	��u��ÈXD���.{+�1�e��l!��>۫��]NA&]����ĝ�ى��?��˶���u��0v{�)��-|��;��dO\>�� ҵ]�ݛ{"�W�CK���K���mP�>�,:�m�(��
?X����� ��2A�Y�{<EP���V�����x)��@�z@/Irs�;�4����D��.M}\�XbTnpS^7���C3$dbZ�������'�)�G�L�o����T�]O��k��-JOܮ(��l�̨NSsz���1`e�f�f�����5+H����\E��y><In��kD1�מ��I�Ψ�J�|ĬcK���fʠ��
|ݣ�Vxh��Z�B��v
�t��J%�k���"����#�əf��y�0�56;���'�M��U�a�P��ݡ����I��?�F�p��)-���8Q�����M��4<C�a���x���9������H��a��NEDߴ3��}���i���A���vK{g"��� D�,�jˑF}Y�2N��Ї�x���GU�w�V^?k���&�a��ѳ]r�e��gW��ܺ�?De�O�/�]��NC�g~��39s���AAm�!^�����v+�t�O������xp{��R��y5���z�h�k�~l 3��~A��Z�z���T"���`y�<G��>����f/\��u����%�&�'�k&��uJW��A���X���0Rr���zޡ�2�9CP���i}�����7Gnkϱ'���8�v4��&���Z�SF�N\�MD����r��������Pp�$�� q�>|ys�����'<kg]f�(W�o#��M���0�m{T�v�Ş�B��7�+(���0SrB���3�K�ؙ��p��U�D��e����+p�Xv-�tU�yǸ����Lo�
�����oi,m�N��G��3��UDR�C&�V�&a���f�Нe��G���̋_C�+�Y�o	Fw�we���L����\GC��:�e�tj>��]'�+h��׏Bo�z�
ۨaI�% �r���q���yR���\�Z�G�{�������l���8�ø�-X�6�FT�)L�x�۝t�'�9��PK�S%�G8 Nv�bMƟ��'_�)D�?o@[nC��
)�L>��;��q$N����6�=9fE��4;��#��X�-;7B#s�f/m�2�-�)e��J{���7�l�=�k7�U�� �2(�e1����?��b�p#��H�N�q�rCrt�f�i�H}N���lƩg��9wg���L0������0�!'F���d)�
!��N��2�~D0����M��8ΰ�7+k,��%��Θи�!���b9����X��k��ێ���p5�tR���� uH��s��,ɻ��r�5��f,��:����S��!
�J1{T����D[�H2�ge��������~7v� ���`�^����������t��V��lF���/ K5$E�g�Hg���
�!?A��,���;E��U�ʍ;�郵�3�5��2�8�e��}��R�C�~�������ý��{�6{�ޤ�D^{---%����YY�Vb����&Ab���Uq,�	�EfN<�pu�֐S����H�@�	q� �D:�0���x_�pAC4�|��ȓ~D�|�n���ö�U�:�f0& T��آ�猻CM6m"�q�\�7O��9�� �B���̖v.�J<�pU�k�d��Ҹܱ���=�d��87��V�.6���sTU��r��=7'���W�x��"d3��:�x�Љ�3�Qt�-���n��He��O��+�M��U0�gU�k���{��ϲ�jeK�GTV�{��� ���s�K>������3&���B^��Q�:�O�s�� ��{sA1���)�aґ�(�5�v'<L:�D?Ӿ2���`uj�V�D�Ɏ?�XQS��w�2�i ���b⥦	����cMQJ�ܬ*��l�g}<�A��n�3(�U�7��(������V{�����E&�G!�V�����c�i�����?:��:�3����r�#B�5ݪu�0F-85��x4q��d�ŕ��:YCx��T�=iC��i�PrɎ\X�5%>?r�J��#r?B*�}z�+��"�*����'��U��p��`�Mh0P�����2���2<(��<�ať����N:�7)���34�0�9�;㭑�����Pܷ��AX`Iϐ�f���ڤ��B%J�h�v8�q��$xW��|�n�D0C��)淟y�,�`s�^�X�N�+6[wF�%���G����>��x�oئ�1)  tn!����ݑ���^I�0U��z�KX`����(�#zWS��H/�"=A�aDZ�_�q��잡����v[��&L�h/��,������������`ٵν^�Q��S��oEVy��_=ׄR�V|�Ca%�GC�@�܉~$U���~1�Q;���L�t�P�����׍��B��J-��������Pk#a@?Y�y +'Hn�^�D�N�nk�GJ�E��߽������k"!?���m#�$;�����ɹ��@�2_����Tn����*]/����S�sL�ʄ/Q�b"fܖIۛ+�WCV\��j�\bWS<��r$�$ʰ�[��x<v�G�?0���=�HI���G�KP������`	D ���,A��ĭ�u�,-�HV-�ԗ'J�Ѵӿ�Mo"�-9������ͤ�Պ7��M�a��Mup]\��k-���K����)�O��@!@z!�N��pBb�\0�|x����J��A^ѯ���oq`���g���}'��ϐƙ���qy4�S��r���0I��C:���p�
4.`�1�0��e0v_f{t��`}�j�;��,�:r5� 	KH�?;��m���[s�y\�-��'J��gc�|��:pR38���]rg��%��
��})��ѣ�ĐuU����H�맃���:�_	P�N1��<�p��(�y(4���f�����=!����p�7=��Ϸ!�)��yiuD�V_^�u�X ���Lu�������P���_Vt�X���df��\�jP\g`LAg*#/�Ȣ���_� �Q\��������w	�����f�xH8j*���h�-�yH>�ט�]_��E�΍��K�-��(���� {���#�ŷJ�d���\�焇�se�[ͲG&҈%�[����&���L=���X}�
���"�l���nk��sKi{�&���~,��D%�7ag��-㲕E)j�=��2-\���`�,�
A���v��96ԏ�=Ӷ�~�L�#O4~�Nj֊#V�P Ar��Ξ/n"��~���V����&��	T��e�3$/@��+����#ŋ���B2��ɮ�k�֞}:H*�����D���~��+�6�#��
J�{G4|#�]Pv����H��k�U���#f:�o�Y+��ˉ�T?���$��6�:=�/y����K�¬��0	-ʖ��F�׉.���t:�pWӿ�b��L��{�WFs1�]��_������h�/��đ�U:�H��{�ݞ� 8�[g80���N��5�7�� ���x���H$g���d�Tӕ�$ՎL((���zo�҈�.��Hss4s2ٌx�����+�|d�D���)N�%)��/f��/ö�2!J��V(vYOڴ��$��u˞�+g�8�,FQ��,=��^O`9A��'�X�3�ajuwcl8�~vs��"WT�3��|��I��@2B[ q�>����� �:+2��?��[�!BM�Ѧ�S	_X�dS ��/NoU֒TY-�5�}���������0���]/�Q^54������*��~��0@�3ɃC���r�jK�>���R��w��\Z��?U�|��lc�v.�TYά���2��8���nu����?.@y���,'�5��%�B�U��V{%N�/���Ш�{a�(��KR��?�NL��'АT��G2���N�n�JW>�91�y 9)��m�nYu8O�9rA�h2��me�bǈQ/�
�f���*���e�om�)f���� u����Ex�*W� |	��s�/���oe5�+����n���~����Ҭ.mlB��K����3�m�H?�3_��]�����="ߋ<{�:)A�z�.�{Ȥ�uр2A_�~�h|04�jø[���r�S��4 K	#������[��S��>�������\$�|-&�h�T���j:D��'n����%�S����.G~�h���5�*��QՋ������f�vn�
")mJv���'/a����(�ƷD��c%� H'w�ӈ�.3����?��[d�;���k��W(�t/��U}&v�%C����WT��v�"I;mYJIw�&��;v�jB��@F����wo�Y�a�'����%�DV�E{��6��B��KM��y�e+�,�d�p��^3�-�V]�G�L��3�W�n'��E�B�O�`��y��ĥ]�p��tMr���X�v-�؋�܊���ˢ���9�� �be��抚zB�R�泃�|��짙Q���N1�*>�^�{s�� ��k�Q'kWN=��.��[��ǎ���<�R��<����F|�̫�~ߝ6ᐓ���H�Zܠ�J�G?\E�6�����`��c���ڒ^T�)��\�w^�(��c[�+� �Z��%n~�/�fh0c�끞 �"<mس*h���'�Z���,؁{QpZ1M}���&z�<��;wlA�������K(P�KR��ҝ�N���F��7�˜�)Sd,�"�T
�ާ	��k�kgj����U�^z�V藎�r�'�Ѽ���US��	��L���B�Ͻ�b�m���SvR���<���z��y���Jə	��4yDx���"��>�S( S����l!�b�gS���ѻ�=��a�Fb�E{��#��V��K�z��7�w�)Z�	q�B�i�h��!�X'���|�Ժ�Vsv[��w�i�zDvD�@�3u�m�2��6ޖ����w��|�H�8@�f/p����2�2�!س��D<标����M�N���9��X������u���@�C�41�Ҕ &c�T���P|�-�]N˵�V8��uZxCi'A�/���'�1�,�WO�EH�\��L�t{���$�<���iTo�X�*�ǹ[�SVR�=`.���z����]���|�Ee�x1�χ�=WP�?�P/P���`
/HK}A�}-L�wi�H�tH��+!��^�Z�Ȗ��4�J���\��=��ln*?�"r�aj����p��|cY�^r�,�����O���W�{�� �
|�~��Ff�%^x��L�r�4r8������s^�>�u�p[�Y�ʍ�k-��\��G��G��}Vg�g�+�V��y{�nl�G)r��ePX�[P��o�|�C�몒av���l�X��'��է,-R�P:O�&�h�Cٰ����P;�i���Y����M}�� 1vނ�p`�X9:|�����d�� 0YD)�/�ֶ�6CNoJA}K�52������.�ycQ��)��3_��/�eb%�'��[R�}��Xs��4��tQ��2�S�b-���C�yq�|?$��<��p���>F�����9�#oAIG��^�4S��&�����1ۋsJnV��us�v)��� Q��g��$�g��t)���T���KG}��@�$��?�H��	N���^������B*H���*<n�p�weI'�����x^H��}�zF���t�:�H��?w^�l�(�?x.�ģЖR[m>c���}�4�y�����|eo��l�ǳG���F��{c&rR��\&�������XP"��L��LS�Xq�L��p��+eΙ���hڡ�]�M�$��w��H�vF2b�:5U�@�%8!')�?z�b��o����ԕ�[��13K--���)��#c��9[��ײ}���������Б���U!�G�(`��~��<,�W��3
���pi�˷�v}D)ju�S�H�:v�ҧD�)'m ��U��-��e�p;��o��[,�<6�F�7$Ċp�;la�6��C�ĺ�Z�9�vW#���4�[��Ҁ�Y�On�����ȥf� ݲaf)���>c�9�.:0X3�'�$���4���&����D�_Z�­�0T�J�+MnL�S � �8�,�r�ז.'�F��ٕA�0Y(�h�Ҧ4��^C�6S@�E�l�>�sQ��r0W��O�N��;7k��
i害z���k�������ٱ�������\7�pG�f/�G��9$��	��{}#ǙK沉��(�l��v�)GL�����b��*�S�������%X��\���Q%56������jM��<]H�_�N�M�20��8��'5�x-�Ǔ��A���IA�,���T��G�(�sAj�uKH�{vKo(޽j7a�B� )�v!�l��a�*�;�bM�� �n*"�"��-b���0yS_�٤yeB��U��ʎ�r��7�0 �����\��J����y�9S��J�|��7]�y\�b"׹�Y��I�[�Y�; �A�T	��J�0}ce�ЛEc��~�Ɩ -�,EL���h��7fǹ���s�d��f�����^���3�k-����Ј(k��SQ+e+��l2+���o�E�#75dJΐ($���1���c���=_HuoS��P`E�@×�ʩ�/��lS�WĒTY^*[��'�Lk��GZ����C�����4�|�y��j���F���Ԑ����{U�Y��?�Xz
(_�<O�`P�)С/�M �|��g%�5Y�)���E.�<RV(6[
�R-N��x������{3���&b�d�-V�%
|;Ⱦh�Y�/�i��aC�A]���J#-��.���Z:��|�n�i�� $m��&���g�vo�Y�9�:cCc�K#�Lk���9�Z*y;:��EB�$`3[����~J���ZSѤ�E�|��g����j�!�0���4q�̳U���c�g�fIk��!T1mGY r"l.Ԯ)%��o�r܄��{vAԡ[�,G!�6�x��bC�*v+:[�Ɩ�c"p����0%q9��" Y��q�\�Æe�t ��C�$7���o��+D�H`�Ԫ�h�84q;��S$�=�%C�:��=Ol��m|A�«R�ڬ*�|���<���6��ˏ["L�����2b;\�+�n:�f�CQ:k`ͻ��wĻ�B,@�_9��r�$j�z�k0��N��x�4^��l���[�	,B��`UFf�� �A��\�0��8�؅3ϼ�<r����e�b֘�jPA�}d���7��B��V�U��k��^_J�W�CTo�ZRN�m������a���I��7����� |)����I�ߏ|qr~5K�P4ws�E���hX5c�L��Q�oGm!+�+Qg��W._�;�ȑ����>�>���:�N�_���JyLD\�;��%*�����xU��2ϋC���'V��6z�twpɣ��o�˘21��ɠ�L�4C� �-�OLXܜ*��#)�!�^�!*�A\����2�¹U9��6]5e.��=(e�N�q�+��u���=lR+�`٪w�E9�ڭ��$��i#�e ^D*�'����m��;w{�N�M������2r�!skHc얐�-��9Y#��0Q5ZT-�-��h��+(��>����� �,]i(Ӗ���D�4m�ҸI��%�l�M��K0A@r&@Ž��y|h�9 �bChU�F�8C\��:r?H~��> A��L��U����q�eA���d�R��	TUxu*<0̋��E]�ft��v=�Jȇ��I�⾭��+
�]liק��H�U���N�l����`C�We�D�N�l�!��c�������y��.`�e���`��4?[vy�D����I}������]��J�lh&7�j�<�Q��K��$lG�����ށLe�1]� �\��T�lĕA]sJS�m�ev���tp2-N���Å{_�`��U��y�N�I(�����:��@c��[���ޙ�l"ԇ��X(��������:tLE�4��-���q��(LGߖ�g|!́TE{7���::���y�&��b�=���h��&����O��~����9t�71�=��^� ���Ӽ�a������$��m�])���MZ��n;�V�؝(ڧ����.wN��$Z�GVz���J� ɮ��q��]�䩗�,�����OᬻfG8�!�RdA���C�p)��"��>�pX��o�P�t��c��OM��v`!y2р��"��a8z���Phj�vU+�&�OM���g����G���E<�׳�����m���PD�5����&�l;9�������,�����H�������Q���P�A8�?RwAzyu.�T��zf�D:-mj���4vx�E�FpV�+A.�)(�Kg�TH�'��x8�I/���u��`Uk��\ߢJ"9�����CX!�Ϯ��ٵ�B��6AN�]�K�#q:��k���+����UN�� �������R S|�g�k���㘦t�z�k��V�xͻ!�8kT�8"�2�ٟ��Kѩ�h�;�l�)��sN�D��x_�>oq�S�";0�a@�A�'��y��W��t�F�.�p\I ���$Pl5��������p#����0*�4 Z���OBд	����	u�Nǧ0t�φ������h��������EH{�rM>׷� 30r_�R�^�cIo�۬��69��.���d�� ��<��S�\s�}��֒ܞ��0�����8̒�4K?��aR�Jf��bS�������n	3�w�v\��Y��^�{Wx2I�*�ɉ���>e!����RU*}!g��*�߽�F���dޘ+��@ͨU��yj�ͥ�Ft��_H��aZ}Z�&�I�=E@�I'��@P����,毕wϛ�`�E�����9+�E}�"_�i���(�	&��7d�y~�C �h�lT0��O2��ނ��a]})#\@/|�9����r�������x��)λ��~�7g��J����2&ɮtÝ�T����Dw���׫,��Ec�!9<�l?��6������`��$�Z���/�����.��;c8i�[ n��J�5����X�Ph�PX�]]�G�s��fY�U�hu���
į�wP��K	��r@[x�r�p�4-�:a���.3�P�^��y�(I�C�WHB��؈��ǘ��Nٿ�:���%�zs�N�Y�^� ) �+�U�#m���@E�o�b��7g�-�J��QS�h�q�\�SJ�p�W���5�_�1jڈ�L�6ot�2_(�7f��� b�(�B�S�DK8�v�ʬ�֨z���=jx=�)������3tr�	yJjΒ;v04:��C1i���4=*z�%��BրE-1�n�d�u�)A��oF@-�^�������Ng��c4{E�o�c�Y]�΅�B��b��&S����N��O?�︨�:�Ё��7��&�CW�acۙ�_s����?�L�-�M��n+�����ě_��4�8��~��Ҫԣ8�J1*A�H�Xba^@�T.��Co|>ta\#N��#��:�"V�V���J$�ʃ�E�8/�[ǋ���R�f����4'����ks��-��h��Ɯr�3dۼ����ӵ�c ���畻��p��{u ;Ċ �_u�R"�Ŧ����9_8���](q��j�B0}D��C�|�Ie��/�LG�v4���;
A�z�1�˟l��ޔ�"�b��c�%���9��/�x��^)�-mkڔ8XY�/?�|΀��,|��
E���j�v�K(�z���߫q:P�N��,
���>R�ڕ����Ң�,����c�����TQ*����w�	���!?��g4b�JBaXZU�	�X�D��%�汖����N�mdN�|�/	F9��ck���8�8�>�1�P��L�HuOw<z9�Z�`��cp0���0r������"C}:�1=�0Q���+)I��A��({�"�t�%R(t&���(.��87�=�.�X"��'f��g}��<GX���1�{��ݲO���0�-	mI.�#�f���47�?���M�2�a�z`C�qH�t�og��S��|�i�xZs���r6 w2Q_�L�gGg������D��IƉA��!�Zl.=dn@��7�c�+�g̿.��I{����)������}6FN���\o����''OG��1V��j�S�3!���Ȃ��^����"pA;��z�ZY��"�ʢp3k���%�4Pr�jb�P�y���̬�����Hm�T�B-@�MC��ֳ�LW����.���Y:>�*Lx�Z6�S���*�N3�v�T��R~RGm���2cE�J_E�YL-�� �g��>j ���\F�Ibe�+�"�c ��_|~��G0R��q��;��d ��R pG�ϻ���g���@�r�8�̮�"MVŹӍ�K�+���S�I��f[�V����[�i���+�*���&3���?��kґO�Mw��Ȣ3	 q�e����|n�r��b�úV�
��U���IY2��'rw�8�`<��_�����|��[��~����7Bo�ᆑ��{�����<��+�<��H���y�ilr�U�S'�-��*�/E͓d./e4:��˲E�h(ud$��Z�&_	�C�I�О�O��1���.��P��	��>�qx�?nY�b�3�R�0�y+������X�aCq���{��� ���N��R��`���9�� ���O� ���X��z��iv|�
�p��0�J77�v���`����%9D7�v��+&�������W���|��+q��Pkӱں��5,��ay��y����ho�^G�O;~i�GZ�`��#j٢nn�בɀ9�<��>J6��\� ��_6���n�5Ě%6�1L�,��I#���D>���a�=�<�����ٱ�?�tUE��Ԉ�(+�*�Y�7����Fe) h�\(,g;^.*ֳ���5�D)ެ���$K�!:S@�]�7��m?�p47�C���QG�w� ���8�_�*��v��E�����	��N��8F&1��ߣ��Q��#��=�A@^7���l�x=�>��?�#k$�bՅF������YC`c*��Y����M�m#إGK_����@�0���%jy'����|3O��5�#f�� �B����Np��X�dC�*��ױ��Wx���!�ۇŢ<������x,	T���D3�O�3M�^�]��}� q0��u���j�0���#�]���f:���W*��;4�ţ��Ё�VP���RE����S!�?�ڴ�Ѵ�yJį�(��U%��j�S=::^�Vm���?��J�5�P���C�S>�D�Qދ�s��#,��-J�4m��=�s�d���J�-@���:�'��}�Arz&���{*���m*6eb@�NP�J�����zrI�|�*L�9��W��;׳�M8|K`8F!uC�+f�ǭL�������͉�b>�@O�^N��	VG�on3���S�0?��)��i�!�O)D�ӷ�&U�]�_Һ���M5[h�M�R��'�=u$����:?���5�'�\{N�y�^/��7x�p����w8��?��w^e���<ӎ�V�k�4d�|I�^��k.�#���m�)��4BW)4�,^gU���~q�~;�O�I���_j.��nl��<:f��Qah��>�l�P{4%NԪb���>��MU�Bgf戼����R�"og���~��jv��٥�L+%� 6�>�I'��z��4El�:n�p��XF�P8��m~����u]t�-�PwLRE�E*��F�F��$o.ə��@��5��b�7�k+�+���x5n#B�v�_rk��]�wX��M��v�0HǬ�����w�C)��@�BK�@Aq���2G�_PZ�Џwȗ�"�e��N�����>7ss�}��>
��_Z��b�ۗ}��A� �S�p�D&��@{�UR��"�}�X�[�/�� }�<)�J�7�j�����2��:*�-������g��Eкd)*)j$���к��M�+;����Ǎ��|���\w��g\��N���*@2���@�>�-��T�F ���a)Q���J�غ��
�z�FWi�F&�J��v�������W����ٳ�6�����M�Am����ţ[�Ul�{Z��d;ex����.����2�ו�c��V:�"UL�M.t�x�uȧ�a_.�%����ʾqa7�L��^ ky��O����I[Kz�4��N̺�_�x�.�Ϗ$�g��i���o+�:��D�$ιI��I�NԽ���z��yR�3j�~��b��wxG���ւw����}��������ܬ�����FJ��;����1۪�_�+9,'��_�m0��2�i�YA�Ir6z:v#DKO9��.Jv:��ZeÏ��u7��n8+6;�����4�G�d�VL��-�d8l܌���������ʌpNT[?�#| D�nƑ����k4a�q1?)�@`�x��t?��>�MPn�L��lX��N&�9�g��IU�������+�	�!�{�z�j^`��3��/�O)�f�����H$����؈%i)�8�'Q�����y7��<������iTd�T��%?j2=�8ts�_b��U g.�	�t���Ș�����Կ��! Ǎ�
�Bw�%�����kea~��\rt )|�˒��=R�FJ�<"�G���5n�z� ��������&5ʫ��f���ZlB�%���qg�+�Kl��_V�*�k����״�&��+J�;h���Dh���v�i�9�6�nYT8}z���i�vVx��U��GP��$yW/�\�c3�z~Ñ���18`�c򞙨'
�Ղ/�n�:�ʹ�|�P�I�<4��̮l���KXء��<���Y����U�N&����/�3�)=�oݝ9�F;U�B5������J�:ڵPG]J�*�:gB�Xe�Yt���8�^���F�D�I���EwS��������+6����o �~�����ӎ�${�O�d�
 g8�%�-ۥ��A�_�.5�(�un+j.xZ��ܠ,���vL��K�
�LӞ��j��-3�&����t�qp[�U �����Z�4"�d�/�*t*�j��^���h�.
����dl�B�4V�6��8���;���>��	0Gu'.�%MǴ��@�o�����E1a��N��T�X=�f�{�L����*R�@�wY�a�_Nv����ۄp�o����"�)�5�ƑF ��1~��HϨ��Ij���k\���bb��:(샣S�=��A�!^�yf��<����%e�ػ�����B���t^.yv�nަ1�pko���9*m?�J2
N"K\�@�w���IL?� C!�;������,�׮��I���@�K��M��7�3��7��Қ��0���G躾�H^���"A�����㪀!Y�1S� �f���O��r���4�&!�E�)�@y�7���×�w��1	����#A;܊����,g�N��ú;O��_���ұ�V�<�U�{�n�ZM�X~��c��Q@[zq�G�mD^飸�]KJn�0}��+Z%�3�ВC�e�Xr���NQ}��^r�N�wO�����4��O	ڣ�\��PP��A�c�ƶ�e�j���MQ��{�^k�/!첺I����pt�U��� .��`!`b���/?JP�ۜ��&6]\V�d���~'CS�C�伸(ts,��x��D�a�N� ,�[F��ў�Tt����Ho}��Y���j&Z"{�W&� xd ��.����Dc���SOc��ac����ЫsW��!��0R=q���
��2zeZ?�z�j�;G�]�?y��*�o5"%���q�hS� 3v&
׶j���>��gI�J{~���P�7�4N���iJ�.��Q3�;�q7�d�oB-�s dP�Wu���"�H4ͭ�FD3�%2U$�(�_4~��b,���2֝`#�p��DIIñ��Y�O��{�L�4����
�aW��}��B^Js���^�1	��֜xű(�?cQ8=�uG�<|�������M�!�Iĩ$�G����:��8�l��&zZ�p|,6��.��s������|譥J�#���@�fIҘ��|��낶��li�'����$ޣ���m�O���E�W�ӗP�,�6(g{��'��$H�ʒ Db}GO;�RQ�m|�������_�Ntq=�>��+CO'Y̰�n�v�θ�~���X@� 0�v3�io��r��f��l�́4�'�Q��lEվOx`�o���RƊ⼹�ke�F�4m�Rj1Ǣ;q%�v#������bPл?�|�U8����������+�,�[�9sZ��O��v��R�C>iBM��^*^;�Ʋ�wմڭ�Қ�����G�R3#��5�4�̨n
Ȼ��������P)Ma_�0|�yH(Y�k�'�6I:�4i�ꎯ�	�=+u>1&f��lL���y�㫨"�̘�,G�2S�+Z��%���J,c
�p��b���m0JX;oyaᰏ� ICs� ��&3��ʄB��Ǜf�l�x��Rj �j)D��:������ôw����	��[��X �O�KT1�J:���}�L�?؅`Jsa��H��P�f
�"}��1Y�
�I^@��U��t{��X���M��k�U]&+$�	��w�Ca�/"⵫+HƵx@�}_�(.S�bN��'��8$��`^��Rh��D$���m�����(5�j����l�4v&M�Phe�U�l^B�n�fC�*è	�CYn�_~�:V2tl�v��������{c �?}����B�kU�/W�A:ꏺ=�⇝=ksdL�繧�V�bR\�����_������4�:������(��6"gj��̐Z��~�cvR;�#7T�e,u`�O�t=:=������'�Lr-��f�z�l�n�C�eh' '3�קP�n��{uW������ICf���[��Ƽ{��O�8?<I~x"i�#���~�-���T�߹��x�2�@�#�1�� ��$�����m�,��و,�
��ʋK�N��q�C�C��� AgK���vX��/8c�6�FY��'�q�t�ߏ�K\���d�o��Ү�ǞJD�S��ˉ|�WJ|+(��Jކ��o��j����ah>�$���ߔx��Ub ��h��L�

+S�r�:kuƱ�L5����G�@�u���+'_[����S� ��qH�'P��ff�4������(q\ê�:�owUJ�}`�7Z��>�C�6j���T������`NX6�$>����\�;�\WAn��{�4#�@9	��R��ޭ��_@���%X��̅�� �U��k��A�l/�?��GhG�@�3h�fǯ�S�t\)A7h����\��;�h	a���u�Y��+����~)!������1�1�I����;T#���y;,��fB���T�e����g�e����;l6�`���3��i����Ь�Y@E/��N�� �ÏLHy0���Xs��-�.��@Ia0���ے
e��0s�9��Z( ��x�'�A���{IZL�n���$�f[.JᑼP ˧���>D�4�O� 9���
�8��_I�g-zx��lN�I�:~W�m��c��g)�LV%�b�;�)�p�T6A���K^��x�J����*��ˁ��a�DY+U]���mn���*�BE�?C"+񗗬��yW�>p,;��H��e�5EC��Eҩj{��>P�:�f�����N�E..R6W�/�k;	o���3!���r�i�v��pE�|�����n�Z��Y 0 �6\ބ��@4����]�+�q���$�t�m1jA�OP?��*��&x��ʔw�	֔������sj���y���	s�n�3�����T���d� �POC<,?����5��>� �*�\ k�[��8U�[4����
���c3xN.�՚p7����#�¥;�'2���t.��X"�!qV���_P%c�I[B��S�h��b;C�2��D��{�FMKu@G�UJ~��=��K�`Ty��X�|3.@Gڬ��-�8D.*��9<���?��"#[%Q(�}��,��q�n��0a�x�KtΘ��m|A�;����Z���[G쪿�ө�>i��)4�՛i�Md-)����l�ޝ$}4�T�3�n:E�o}���Mw����E�sH3@�z[~g�#l#�N�n�(ok�<=T�A��%��h�#Bc`ig~��U�]��HMh��L��Ul0���ѳE��`�r��'>��[�%��M�G9�վe^NvJR��|T.jt�v�D�~P$��P�	Ꝕ��;@���O��������'{m�;��2�"��,,0��u0���o_0��j}o�`�Ķ�m�H"���3��7i)��xhR� C��
�{)0ٯ��_�Qڲ�1�̌'( Z��17���+@�n��@s�;��q���u'��ڔZ$f�ˠ�鈣M��ʉ���#,�PU�j��e����g��y~�G��'װ` ����!��.Ѽ0A&���og"M���-�wO�O
&w)�y�
u�G�.oGэ�-��d4A̧d���q�b@�*o�p8�!5��v�KhfBՏ'��?��T�ؗMX@I?�mU���9���N�)�����M�����������|��L�����e�=�O3z������«e`�>#�?����i?b} ���U(+ئ���:a�J�n\r�����R0���z�����+ؔf,G��սl=��A�D뉎�rWtc�kh	 [�b��%绒AtG*fBϝ�6��7Y!�*������-HK��GT����uh"�3�S��q��Rկ�u^ߪS��C�H\�6u��:@�f
��f�U���ʳp�q �΋4Z��y�l�J/Lb�9� U~��Ω�.��*v� ����7�uWn7��y;�b�ni?�������>����Bk��P�-^��7��a�$�U��H8������=*�S��g|����o��o/({w�ۚ9<y-jP<ȫ��\]Gi��ը�R̰T%�:e����(�6@0��6�G��a1��n��T�@}��=ŵ/��[rآ��=��� &P�v�V��ij�.HH��g�T�m. CPs_{>�Y��^��V����]:�ϳ�p�7��eˠ���nL����1C91��X�Ο���M��a3.#o�/�+��Mb�M���;X�� ��u'��� �k���$��+؟a)lH��#��zc̀�4r�1�%}�5��T������g`���رW;�fW��PR��M��[>n`�\^�N�- �V8JH�F
�?�,`�=JSB��^}�h��h������?��]f�w���CW3�.�3��9|zM�9:��D�\�Qd�����;�X�f@`>8o��X@C�E��X
��u�m%�v�7�^���eEC)p�{޺lh�	q���a¼{L�ø��#�ާ??��e��^�v8=/"����!��{"��4�(���Xv�a?1H�����ۛ)$��4YT�o5�2����S*��D�`�(��<<��ٖ�
&�]*�����E�r���a��}��E�t6k�E�� Me^��'�ƿl��⡴�TO�~��{�q��W2�o�pkO)cΩYR�0H}�#/+�
�VΧV_t�K�a��'F��.�Ӈ�S��8��Z�	M"j8�W�M�����c����rE)%#HX�+���f�6xg�*R�L�fH�,gn<c�4�Γ�A�a��G�P���pP�t��G�����[�Ԓ�l�×?{��B�5޵u0��H�o�ob��J~�˥w,��%%Ч��usF�1@0�c�%�|t��;��'��N�w�5�ף���r/c���Έ=q��YU���vd�[j>��*�_�����;_�\cNR�i#˾>���,Ȋ�We�[p�i�"[�Yh�S�-��$��#pg�Fx�m-�Z�Ví�u4Ym��9tY�NI���\������*�ڽv��[Q���&���F؈?�:}���#i���y�@�=dO�`���K�� PT���V�2A�kf��`��_PEi�~�T��8�.�K�G��WR~[sM�xU��-Q�ӴX��O�'Xn��[�z~��!Ú�m�-�jN��V �a�d�SH֩c�M>�BD�5g8I�l�>� jZ�~�]؞�$J��q[���>�:9��gN��F�h��+�%��'������_�n�c�|IEK�aO/�_4w�_.����ULM��-|�*��ru٧�s���+�~���ר;�I��X"�x�t���T�L�RT�5~�е��ɟ�2��ogM��	��NhJM�uo�M�,��d}��W�D�"8��w�
���Dd��.8���v�OF���%���:G��(�t�� L	"��Ylf��*�ͽ�H���"��]�1����ӚS��t���[N���&߈7�Ȝ�Z�PF��Bb�Jd��:�fE��x������<��1��4�I�2���QC��B9V3s���.���3�����U�mw�*�!v%�g~0�fDw�h38L�S3��{��1d*$�TXCX���9�|�k"89:��m�b��^�0��,&��͆Y�s�G���z��r��j����2-�� ׃�[\�I`�\�?�=���y�Og#��ƈ��[4�S�Ñ�=t>N{���g�'�3�GL���L��į0�h��>�?Ҹ���1(!��Q<BɆo_R����`��ۣ|R��n5Wߔ5>���	�rC��2��;�'a��J<�����	h�oj��B�~��T�>���\���װ�(��g4�<����m~��C���t���z��!��4�%��p���[Է1Da���(��ftҎU�K�d�?\�)�m��s��|7��x1hK���8h����D	��m -U9)����LȴqBwo֌bne-����1���Vܞ�6� ຩ,h���Vx(#�4]c����h�Mh�O˦��W��l��l<�����Dj����rz<|E����ы"A�s�Pt!1!�j�SԆ�׌? Ŧ�l���1�����xQ���~aO(N��u�G��t��%Ԭ�Ŋgwh�T���Rl�Gg#֝�B؊dNO���W��Z+�o�j|�I��ҥ�m�M�d�2v��Eڲl���+_VP_�V����;�S��c�S��W����7�'<��ŽS���Jg�5@��~����21A��1Txӥ�cE���x���EB����!��`o7f�����{;0	���!��"�t�r�lR% �l�����k�b-}���-�M�h�8`�%[��d8<��g�DD�/��}�8�}n;NS1�b���^P'[����
τ�&��iX$c��_�hJ�N�}ÿ��>�cL�g�����{w��J ���}�Z,��EU7�{� H��.����nV�$X?�&��pb�/�7�$��H?׉Ŭ�6��ȓBq��Э9*HI�&�-=���rA�\ń-6����ºm��1r�&��4�\��bg��p!\���g�	TX�҂_���.c�(V�:�"x�݂8�W(�&���ƨWI�v5�qל͡����1G��o�U�K#M�@'>�G��~H6�`-0Oe�{8`Y�S�2�dAۻ��}c�5]�D�g����(z��B����2R�X�$��Q���D�1��0('�t_��4�����J2��
ŪB~��Y
Vy��_�^q���ʥ�>�(ގ�5�uv`��h@�ut�c� ��0Ou:l���lo*�p�clx��#�e���p�!�a����w��.<9����K�8�Z�q&�nC,�Jh,�S�hUkE9�~b��[�P"��2l�}>8[�Y��X-BG#�6���X����\��ú��[e����k���-h�4�+�hK5�]�M�ܟ�����Ww�I��tP�|Q�������`���� �$:ӣ���=�,'�A���1�$������)x�P�Z^���-¢8�k��3H�HN��fA����z̸����W��D:S�M˕��3NB۾�F�=ƛY&��I���<��^�-�5`B�P��Ro�.`��
���whh�1ā��B�@�~ՅG�qF��OeTٸn�h)��샐��8�-�����9v���1�9	v�{��R�D�Ve�77yu}��GR�̅p��TR����K���IB���}j�.��3�����#O�@��s���.�����B*�m�h*��g�}����v���:�,���w��'������j����
�7�7@�D�>
Թ�Ԓ�%-������i탍��}���+�5���1n�}#�tӟp.5`䍜Z���Q�ޓݙ��g�@QYqXxD*]��uf3ك!n�ѵ���H��\��[�?�M��@$��l#j����m���4RD}��n5Q��HzM~��=���u��@n��<_���زr�8����=�ъ��0Cv� K�ca9�կ�É�Wx�����r
�服�5�
߻
"�g��B ��_�sμ�N0��[�h?ݍW���\F��(�E�S{�Lѻ>ӛf�(3bo�*����F+p�{�N�3��B�ي'iXmK&������O��T� �nO�i�� ��ׯ]� � fSz�n��,,��V���=�u;-��:Y
.��t:j�� �C�]?��IZ�FN$S¯.�a;���hUĽ�^
cO[4K*��8ُ�G��� T���Z�>J��z`�p��3atpkL}�<bE���"㒀A�2Tg�I3��x�2+�^ ���FD��v����n���{|iL0�朙ܾ��X^qB,���H����Q$ b�e���rf�tc���A���S
�w�O@p�c�Y���v�HU���M/��:��17'�}D��P��G�j�7o�� V�3�e,#ie[��e��=+�Swމ��W#������[Ӹϸ���D̓��˶�uş�j��M%U��S�)��E��a��73�ym`*(�o|���<�8J�k"�������u��.-#���2�� #_��q�$�-��W�w�"���*P ���"�o3j�7��>4A�giR�j/�� ��&i�L�li��~uI� ZiZI��R��l'f�FHo�v���#MC�}F������:��gKG����H>�l���1��X�E�JEl�&+���b��t�r��)B�h�㾚�����62�� �Q�f�	(�M���ƀw�j��g*�����CC�mp�YN\߱2l�=j��PD�g�g�x��UE.ƈ�>��Xqv��|�;�.[�{f� �u�@5�N&���ىua�n���H��\���,e��Þd9�Ò:3�AޒF5�ݨi��`�Nh5�p��v������;4�V�5��uOD@|�@i�l��j+��.��p��$t�&�d�Ҁ������+�y �����U�$��5���K$E%��)�GӒѸ�l�K�"�$��"(�_i���%�{?|���+,��_�� ߰>`ޞ���P6�H�osX���Xp��dS3�?�_s�p�t�XMàڟ��[�u��GǹN-ؚ)7ē�ݺ���#�A�����&t���{e�y끯�Ve�;��}����5��F~���z��NS�	����ԭ�:�o7�+����4�wv�t�H�Xؾ�J����SB| �u����@��ȎRe���%�2"�_.'ъ�Yэ���1x*ZEB��'��M*���'Ⱥ�_?\LZ�@q6�����;�k
��As/#V�[,[�2(�T���Ƒx��R��^�;�qL�,��5qE���Qo�����ǠӗXả��uku�Fݻ#K�Q�9�M�N�:�p+u�n�z��ݶ���b+���+	S2 �����6�YS��N%�^�i�O�^����ω&����5��^�@j" ��tJ��l({����6�%4���V���F�D�6i�P�'���'���eE�L��|>�-�o�]��ohv�˥�nᕑg8)�ƣ1:�N����JJ�<��)иW�*�w�(�ֵ��f�����q�r/�L�<�7Y7�΅b&���Yx���oG7~�S6<e���n49*a�PbQ+
ۨ�����?�1R?x�o�����D�S9[�N��l߶}H�R�^��~_�Ә6�j�l+	X�"����A��+���� �Ǩ�)F�ǋ����]��F������_�%u.�~QH�=���@� � ���I�y��I�b�]�����v5?
�{P���Dh@rII=�/&�p�/��m+�*Ԇ��n�@AS����D�U�5�ݮt��r~�$���p(�I����gp�l����RW����B[[|��q�@������D�2�bs�i)��!dv���z�@��#�9 ��X�1���3��Rt�����H�V[�����,U/�/�����5%
�LBuhВ%��JXK��-/gۢ���qʪ�����!%pf��2�0��0�"�w(���)δ�B}�vߋ�;5Ϣ��Ω�i#�r�F=M��}�I~W{k������ݰ>3�QQF�|Qs���=yH��͙`�L�a����,��� 9���~����:*Ny�弦[)�C%�o�mM1��� �4�v�9��(7T��F>��)�Z�_�&: ��r���#0 3��g�����uP��e]�K~�3����-��"���o�)q�|��ρ���s1�n���`�ο$�x��}���8s
�_\�/�hj"B��W�"Sj�yZ�����?p�Uw&p"��|���ӹK/	ɹ�+��}i����{��b3)1sH"�FKh��v�'J�hj�@���Ie������*��&k��js_��~�_?����8%�g�m⾉�Wf�$�T2�們�v[���}}�g!x���މ̔[�s�vZU�xY�.!lY��x�]���v��s�vF��Q�L(�W�x�TN��<�W��2���[4������#e���6J!W��R(��� FHb-�0�!3Ғ���wr[F�~u.AU����,,0h{"���b��.��0�Qaei���"tHH��k�o����� W�+��h�O�_X�D�w�ɜDW>��p���ޙE칈2CT�^QF����u��N��BRZ�7�lI=�q��er��췷��A9�|��Z���*�G?������.�����1w�y�&�}�I�4�����F�C�'Y�l��N�;�R����'Y�?����_�X�e���[�&��`��pJ	�`1c�����)ψHV�������1+���;�@Y3�Sz")�8��Q�x����Gf�ċ8=l[�]�]�o���1�N��j?>�l���)0��c�Uo5e�{ ϓ=�Q��A�Rn]�	;P�nO.΅hB�vrQ"�c?V��PSOK�jB��;'k%�� .����6����#�gC#G0 ��t'��T�1�
@��o%�l;�ڔ����
���7t���_"����a������T�&$F��.��4��5�f&7W ��F ѡ��*�i|xcq�W�����n� 8�2�%�o�[�6�[����VjLƇnk�amjb�pZ?�ɞ�06��O������G�"juX�e~�QǦ�M�c���_7�y{{��SmՐ���Y%=H��^���i�q����]Uq.�Z'0b�R�I�ŗ��>H���>[�m 3-�{r<��tV �#��Hԝ	bh@�u�CS�����ǐ�G<AV��MaB���n�J�����+G�T�=�ßBl:�����W��Vͯ��5&�e�3�kH��Ϗ~O?��l~c�|AY�����%8+0�@�l��T���$A�?o�a٪���~Ÿ%//}rw~��;��"���N�&�1f=ZH\e"������l �9�Qϕ�3��*,@�c��3�e�]�M�e�q,	E�ox��j{����?���(��l�~1t��	�͑�܏��r���d�H��!�[ l�vӴ��)�]��U)R��1��ưDԅ��s�N�Bo�x:�NX�JN���ƮfnN�����ng���M�0�^H�o�n�!�*-
.o�� ��,"��g�khF/�'��J�`��YN����B�H���0}eo���̷��w:��g��ꅼK�<�f
���!/�26N,2��A�<7i�˛�~�Sw۾��$�ؔ��b7�Y��m��{�|^B���-1���^��w��!az�l���΄Zo�z�,������g}�X�}��-s�Pd��n���$�)�y(������9�3��xe!�>�&�p���A�o�\>�RB��8�a�:$4��m�).��4��sE됝a]t�����u �=�z�� k�����|@$�w�U[�hҩ�oW�A��*�C~���E��I��pm��;�h�I�����Rx�J��ꪜ������|�~�N6�t�y|�K�h�O��"�>s�c�G�R�#��ju+wQ��]�i��M���{�\؆�Zi{f��r��''�߅@�{�F�W*SU^��%2���0�'�\�e�dZT��^�8��9f�!I$GS�u�f�<�u�}����_��wX��Yq�5�?���
����zs����hU�`\2ON/�T_+�e_��Y2!�2��\�����H�8���>�B����oh�Q���?뙷q�=9��G9���e/��@�n��p�Pg��2�=�*p)�e�H�<��\��/�j���B��s+Z��>v����hw;,���=��d+7�{�)�]�7��	`��VЫ��r�
��6"�� �pqL�#�fdF"á��uw��G��}0�%����:Y�$�4�4��!��<� ̌AdSBvİĳ(�v�܈Ǣա�f6�O:Z�����$N&��Q��p��W����(���q�
��Z��D�7U	xc���$�1�`qIV�)80�J�&�+}�����ށ��B�� �^�Y»\�׈�lS��2�<QR_'[
��V�g��r>o�^�B�^ׁ&�}��mDPa��;�CިpL�����K�V� 5���A�dH=U���C������J��½�^��ԗ� p��$��t�@M��[����Ǐu�)����޶3�%V�K5|��Pm8}XAd �1�
��{ŝ�Q���Ŧi��l�L8��X
A+c"�$�a���3��Knk�X�����[�df.��ĩ��oXiVN"�1o"(`/�X����.ӽx:�g�V���x����"�t��=4�-#4d!�*$x�i6\�A{�,GI��^��@�0]Oy�9�����h�C�Uk�VU�aM��6�Q������@g�.͂e�r�C놼�`��&�c������u.9��9 g�rh�o;r���Ai;�<&���ߚw#��<�F�9��5���p(���D�0�t��~LUܬW�j�c�~�Ĵ�	�������bz��Ο�J,D�[KnÌ��z��tj�5�#��_��];J�2���M.`��)U��R\�[�Z!�M;8O������3��n:���<�P'|�<�VAX�����c���y6�m�/6�:�c4��3�V�9ǫ���!��6X�_�~���T捭�*!xc�	HX��i�7Q�S��z;���]P6iK�g�n>����ɖ���f�!g��}L�d*�U�ӈX�Ϝ��q��m5}wiGM�MUR快Ä����EB5i��US��6+��i1��6+X#^�4�������6}W�Q��[���h)q��6��
(��^]#�oK	J����%8��5�zq��4�^N�߂�kC�GX�|U�ƅф����D���Э婍�=��œ�)�%���Đ�#"~j�E����*�Sٶ�oZ���j~zA�3Y�A���V�[-4 wdd���aYGSĔP����^-�R�1�aj�@������d@DUx�ٺ�����7b���h%5߆�ڈ^`Y����|��S@�,������_򅩀 Բ�w����Ęן��y(u�*o�9@jr!4"�ࡷ���ۅ��a�Η��4S��l]}��F-���58,��$~ͫ���O/��0v��Q�t���p��ū�G���02b*g��q��۫-�vL�9U���Z�/�P��@�� =rEl;��q81#?���/�8eM�,��de<b~��@JZl,&�V�^�(߀�.������7��I�]�;d ��ݔ.�t�  L�7v���}�6�2q�gXdPB4�nw�,�hq��=wk>!�k�a��aAN���]UR���Wm]?[ ���@6��%��L��Ur��P�3�]�&�MA�Z�yF�d-2;�<�X��Pu�҄�RW�j`,h9YL�2��ӄ�l��w�q`n�L�9�E�Ys�4O�)&���ߘPN��0|���߱9̋h!��T:����Fi����b�e�0�}߰w��]��+64��5K;׃��}r�-P��_G��:b�-�/�vT-���#?P$^���oQL�Ty*�uY��	a�r�Q
,,����zY��_��S�ծ�ʇS�%��0���U���I�e@��X�OCW)B@��׹H��P;a��-�qFu�0�6�u�����[���CH���Ud��3KO��x\����6�oU�D�T�P0��ޒ��|7�޳iII�j�##�L땩�[y2yiN�ՅXz�!8C�q��&=8Q���ѫ�%��OD�C�ԝ��.�q34LƁJI�Q�(K�5���\>�J�,hQ�Z���t�y��tE���U�A�̫�z��F���HJ�]�>���1&Ґi��EWM.T�>��+�(��<���؃�gԸ�X��c�DP����=�eg�{�Nt��;� ����YOjSY��q �Qq�{Ie-_^�G&T��q8 ��t���z+U���p�`,�����˓wT�I��F�v0UXp����
�|6ɓD�9A�/P�a�	��1�ͮ2hT���l OY�T��9��+4����d|��BD��uΡR:�����1�x:��;4����� �OS�U�
} ���#�O�󻡯�'���_9���J���F���@�Y1��wEQ*�+�Yd����AI�r'��>4˿o���Gji������z��
l�7H_,J�i�#��h�!@*y�$4�5ޕq����Ԓ�T�qz��,�|���'ٟl����4V�z�F���Ncl[��޵L�	���s�f�o��w ��y!#X�����g H{|Iș3'��*�∬j #�i���
�|��BI���-u�|���߭��+��naͿ}�>Z�a�0�Ku�ge�NJ  �t��u�>I�*{����ZA����M��N\�s��,Yy.�>T"�%[C���������ascV�������4Trm�E�B���}(Q�T��V��)�̪N������J�iET�qOeh~�X� w�6V�^ȫI7�'�7.tr�����y��k��u��Y�T2���0���^oNd9�0c<�ab���F�>����6���]��9��~��Ή�1}ܻ��O[d�_� �Fec"��9%�
������3OwD_E1H>�w�n�L�y�GT����Y�=�9�T���,�����%�nx�:i���mD���h>���doՉ8�h�\��`�A�&\�.�`J+B�ܘ�	�Y�R6-M�j��*�z/+�3V��i���w�Y����q]G=yr^mF�R��%�l�A4@j<1���{w� �Rv�祢�����
�\�?9�8��p�zҿ�"�=͂������h�z1u�cj͕�;Nk,ۏ��,���w!��$����}��-L04:�Ɲ'o�n��m�uF�V�[���"������k�VT2c��ФP	���/y7���,��Ӧ���z~��q8[��`{lӤ����	�f��ZtZSܗc�j7o$�y���P��FLG���Y���r���֐m������)+�.	��)��!-K��I�����)�T���]�-�x]9��$ �����k?�Y��Z�פO�8C�0�N�3����˲�mT-7���pd"��3Ћ~ݠ% ���G�߯_�ӗ��'8��e;^�J����p����{�*OUrKc#�:$�0�L9��4ȍԲ*���|w%c�i��R/�0��6�|B�p��bU��S�2D�ZMg�z�]��ǭ�'@D�B� �p�;� �{�ي��U�&��^��iV��Td!�~�r������nЬ\{0n��+v2�I��ܾ�Y2�J�'y�ӂD.����I�sb�[֏�qK~�]#�D�d�6?1�}
����ث��]�M�~ )�����kJ���y?d�ߐzG�r7e5��?�{�X�-_�kK�gB-c`��mM�%9�����m���[�틥�����$�W�Z/�3?u��LPV��^E��jWk"�r�����+��gB�P�.�\�2\�Z-"Ҫo\"K��_uW��z��/�Ѿ���fv�KL?m�)�O�UP(�^��?�S��~īM8�Q�dm�M	�+�h�NW��L����1��rYQ�+��[�4_�x	� 5@.�q�g����D�,�!�h��~��������a��h��\���#�vjÞ�����qT\�V�����Y���)�n�l��c�ȁ7 �y�����x>�C�d��Ƈ����BL����k��ѿ5�7v���?H��o�	�����&va�ܒ<XqT�:��W/yKf������rjɫ��8�/ƿ��un�����M����	�� Ӗ�(%}����;e�\Gf;Z�u+�i
�r[L�M�t�����`�-��X��i,5Yh�VKCM%��,��r� �x#�w�tE%{�f�i�:Z��$��.��d��h�� [d.��ٔ��������#�����6�b5��=��錬�q(���]��/^�;-
]{#�9��%��0�:޼�@��]��-��h���W�ߴ�g`8�@�)�%�s1cFPu6�ؼ���->|�LT��?�o����v��P����-r!����@mM�qQ��]�(/	�)��y�-epd�f��W_�u���g��k��k!�o1�,X6��F��#Jz�������g�偸*=�����\��3��X�d�jX�Ƨj��M�z'⽠$�ѩR�m�fc=�c����EB�c�r��ycg-YT�`s�\}���R0���{�h���U ?��EL�n�v��kd�y��g��d�&��!R�L�B��ƀ���\�H��30#h�jI2�N�W	�s�&**�W�F=�<���T�å�b@J����~���4�w�8�Oi�5�n,�2�nB�l�:���{��ْ�R��G�;��q).q���tT�S�v� eQ뮝{�����;r�Ck4*2sP���S���S���7���#_+*/���cC�:g,�^j��AmU�S�䐜��gL�����R�J�����y'�/�I��&y&1S�5�����ΎlN���+g�W�m�ӫ_.<� aC��LPI;� v��HB����o,r�`݄2h�,�M�����}<��n��/I%9KOI-s�f%D�ƈ
jI/U��є��8��my��<�t{ko�У����R�
�g�@�T���Î롴��HLM~j�@����3�3��M�!���k�u�O�`��
�/7��9�&[�0>}S��#�7j#��x����\��t�lI�'i�86L�;�(ucA�ns�����DZ#��:	�'��9�$�Sl
�P*���m�#B�����_�F�C wXm�"�U�g�7�7�ߨ#�훨�,���Qޟs_?��i���>b�-O4$�埜�Xm*30�xx�46q��R�^öa�^����O�	����l�Gv;]Ak`������F�J�����w2�n4��ĸ��&)O{�iŮ1r5��f�ŭB��\�t��U�{�$������W��͟P��T�t>v�M��շ98<��_�
U�ˤu[lˇEw�F��Ke|f�L�f���,:��W����'o�����uT��w��x� 惶�#m�S����'"�eV�o�t��Z�I�E,�>�,s,�*�S��P��l�N@�S�b�p�?���	�Q�_�����H���
y�=xR8(:D�����n���y��+\̫���H�ϗ���7���ܽhk�ci⧤l|A�f����%�3pYԅ�����âW&�m>�5~�G�
't(`�>�gT��c��G/���,(mч��ܾ�G�.c�@�eq�m�V{��cj�$�A�q#���Xcy;ᓼ�tǴ�=���|�=4	N֦_�E��7A�!H*ɶ|��ccmƎ�}UA����R��U|�T��m5X�F�w��}�d���RF9s���Մ8�
�$�V�"h�w oBp ̷�m�Q��u�������N�6����P�>��s�cKV�QL�J�JNEؾ�`�F��J��]^�k���Gn*�!��л�� Wo�
S��o ��B������ݪB��!��m.Q��᤿��q�s2��!����\tr��2 �E��gSO��}��  䫶�aY�`�W��_�l?j��+��R��(��<I�r��t���9���,۲������a���:������m�"@������U��rq�W!�y�(k�}���Z�]o��ƝsT�%X̞�O���ű%��l�t�U�d�}F�6���g��I�q�[����=����	��}�mӚ[0���б�/�[i����đ�z�$��R�����QX�ws����^�5����K�V��l�^�_}w����H	5�"�� �o���*�| (T�>�s��Y�T�H�u��$��� x�'��ު}p�9p��>{�h�.�`��>{�e<N�Z����Z��o�!n�z�fIH{�7g&�`��>�}L������B��>�U�G�|�~㮺ǅ*_��DLL��
�*(k�cR~cPgN��|M�x|A�����4��ݒl���g��L�Ȃ���(�m���у�IO��'9��,R��B2�ʜ��"�K+�E$ǐ���ϑ��O鮲�	5Y��u{�W�B�5W_��	�o��z��;m�{Q�E7@5������n�_0|�#~5����a&Ѓ�t:��5r��lQ1G��N�"���Ǵ�:�y������` �{�ߵ0-]6E?�o3I��U�	qX�]xf�6�eW&���Lg�@4�*�K6�3Ր�&^|���a)�^M_,�fq%z�;P>�gq��u���T�J������k�K�2��l���v��
�kW��0�-���.''t!���0[���x���VM�ۻ�b�����l�3Y0����A���� ]2���d`�]:w��Y�flS��nS
�	��1�����3���,��g�au��ۮf3c���r]�y�g��ĉ�Z�#�������pI&W(ɭ�_$�4:Y�$����K�".AUx�=2�ϭ��m��mS���4�&V��*L�$/�CYbi��-�B�4p7%Y��(���ǩ��,s����[�m�9�q�}����!��y�I+�w� � N9]�Y���=�F�)§D�zs��N�s�GX��B���Erhە%�-�t�]<��%|TF^�>��r��%��2{� ?X����˯�K���YVʪ�Lz�U���N�ƀ����Q��*��6�i��$:�֬����o���� `�&PM���:	�gid�p�S�0��"�ђ��c���əN��Y<����<�h����R�w�/�@�m�E�Q�tA���Ἁ���������mT6��&̫G���Q�ZB)�*[g���׻B�J�� ��Y>��w���A�c�h#`�W�(���n�Qn�#��}3�u�v�]�q�s�k*�c�N�4XϪ���*5�D�B�y�������<]xu��
J���̻��]i���%��-�6P��Ԁ�2{��.�	B֣�-_��n��w"����x�aX_,�]'�v��X��ߞ��N��-PF��Ci��ӝ�������;������)τ�	ˈH� e4�x���ǜ��n���h�o���J
ԃ^0��E��f�wkk��"5h�ړ�Fe��UCC7�W�4���_�i(��hD<'��&����̼�uf�������荄��*2�A�jI�5��zN-���B7U?�S6���Z�R�)nu{�~w���JO�'G����)�1�S:e��=|
u�QP����i�N��Y��i��I�ʂR�ٞ���X=���7[�^T.kU@�e�(}�u<�m8��l\�v^s�e-��\�Gn|����h7؇��DC�M#���ȇmp%��US�,b�!C�~Ԃ� 1&�K(��OIa�jc��<��x���'���h���l����Tt��fn�b�	ƈ��1T�.��	���I�u~�?sZS�Ԃ)n�����s@��N��9�����i�څȺj�	��Q'�m�tr_j�L�+�Q���D1��������B�I���w��/3�G䦣E�
�B4���Q;�9��Y�c��K�T<�4!R��y��~���OH~�/ވzStc������1t�A�}�N����{�:��%�I|"XvZ����h׭�]�1~��fK=���GS����"]:T�! �8qK�»5+�%�����#�j�� }����o�,�e��O]4�ﮈ��fwټj��,_�����+��I^#�Ǯ�ӑ�9&����f��nr�4H��h����)��_�z�C��W_GH�	C�Y5a�>(����pk�,�}䴠�j<�D�Y�CfI#A���T4S�:$�;���sm�WGe�"��Q�`�va�t4�S��)��U;�؊�@�K�E����r�	�kc����J�K�����W�v���t��<9jq�%�-cv��r(㇁?���n���2�8>I�F����X�6q}ϲ��i�wi�h���geP��d�F?�����ł��{���k�q-	j(�����u�Y5$E����۰�D��G �HVSm�N����[rA{	l|7�4��|X�u�9���{���f��&`LZCs.{ �kI����j����8�}�qj�*�G��d�Ҕ���\!�J&�;�[A�B�j�<#?p?K%G\0�:Ȟ��hc�"�â����mf�Ц�=@���`Ѿ�Y�2Y�W��9\wI�;�3)p
Y4��ʠ���!=yu7��-gH�m���a�	�F�����%Nӧ��8�w��J��2���
��rg��w8�Xf���k>�^�2�ZZD�k�8>�D�}�֊$L`��h�K�5��À����cݫt����4|�ל��+���pM�~�T��=V��sgD;	���!�[̸�tk�;D+�p�ʯ�-y�t��o,=|��S�\&W���h���{�GM��:4�\��is�X��Y�d��� �T_o�C�tw6G0c֠{QK^�m%��*�Կ�ve�D��j��+bw���T���������-n�m��|>��s�5^-h(3C��x[�i�8p�v�%��ˆҎc��~T
XG4�<�y�5{<��^��i�\c��ڹ��bY\_��-_Yc1k@���2bk��k�u�#�����A!K�%�����PS���G���^�{�RL��G�����Jؙa;������Q&Y�b���z?:��n�
b]�M��M�:�Eʂ��ȗ���,&��C��[����;��aIQ"���#��HR�/z �x�2�@?Zzx��K!�(�y����AD�>��z��ި���R,��$�Y% {�Po�O�1�����p�彂��c'�!���v��M��X���M,���S32�H�e�,���ۺ������S�p�I���������m߀���>y��B0�6xij��D�j�h�+���ҕ46|;�W����}S0�������5�t�6���aː�:kk�`B^�&��e%p�v����@f�3�Vw�o��m���f�Z<�b�%Qv^�(�.��l����2�x��޽�3����-kH�����
]=�S���C�u�*�e��xҊ����B��(�-(Ye��:CK�4�Q+TYE���~kGIA� !δd�4��� �/���� �޽r�Op�)����Y^�8�=�]�`�4r�P����cf�Jyg߅���DS��y�y��!��r+	e)^7ї	�t�{K��%�T��oOa�P�U++z�!FHQ�gL�Bj�����qj5����v���H`�����#�#-�]�}kLl+����(E��Q,]r�b{�1�FD�#�
N���s�ז��df	��}=0o�~J���ffd%���԰i5�ZK�߉p��vU��C�iC���]��r&h��=F�9R��f��F\	R��@��AL5.v2�������8��!���j� ���8<e�������=����V��߮_o�]����Z\�:]Sm�V#��PVRaq���q�h}>�q�wR_���P�����R��!�Z��I�ʸ7{�o� ����=��7�8t�!q��A#	�@'�\�""��"�߻�/����[�p�����3�'�(��gRO�kx1pB/	�<�*�ו��6P�"�u�>D��QA=�i�"F���C��K �/�F��ַ2����e��͡*ek�x�|���3�c��b�
uv_Yĩ8�P.6�P��ڄ�#�t�#}#&1�+sg�����^ö �]�(��	\�C��bw
/b7�,�G�
��5�
�k��D��O�X�T<�n�
忥)�9�馊zQ��">�̡̌��?zu���zA����ś�����o wR8	�� Ͳ];Q��pTd퓸��Iq�J�(��3ը����{xvNy�(����=e[o
хb�px�W�~�{#+۱ީ����w�Bm��j��)�T����52o�a�N��f$���UO��6���E]�Y��p������/���b���b�3��l��ÂZ��2�<��������k]ś���|HF��]��
�7�K�%�����N=���� ��Iʑ_�l6H�bOa��,AI�$�+�e������$����r^z/?�i�Њ%�0x�*m�U�h�4Pk&Ɔ�X����>�y=&��y� (�Hn�$���\��R`̨��y�>\���[���ĭ�_$�q�-�-ɕ��#H`>��SJ�T>�{�ö́1��>��4�fn-Sȓ�QȒ��p}akg�)�/ʸҐGH��5+�nQ�c�7G�g��~��ޜ�f������Х��~j!U���Q����	^0��p�A�BC��D-���~����Z�E`����q5�k�j��������qEZ^�N(�XEϓ4���m�	��n<ݾ�4��"x��C��b Ǽ�@���6{�����;�@4�z��㬖��X�q���������V���D���i�>����9�?�	1�C�>��9"I&2���i�W6�EF��`iQ]��-���{���S̅0JB4�J'`�h�y^ߧ�"ù>�Ae�y')�� ����;%����L�5~=� H��2c6�2�;�5��r�2�Ff�)G����eMIM�m�-�Q|ܘ!p���|�D���&.Z�l/{Ly Kj2����Q���g(tjO�|��F�T�x���;"$.�-a��	n�Q3^�����F�c�L�d�9'���}6�E���SL�d������pV{�t��v�kk����8�>�ݾƆ���_�-@B�T�$�}S��N��ݫ�;`��)uJ^��{�#�	p�r��fK~�����t�l�����ﹷ�D�C�;c�i<����w����둭�R�J
�d�Թ誽Уkounh��J�@��JA%��J�X��P�}�5��_:���Y����^��`�3d�cX弎V�s �,z�F�u��2�@Z�£�ȍ��e>��ne�%���IB+� ,���)��b�:LQ�1�����_BB"�
��N!�B�X5��sK���䋃A	�g@��^�N$߆�䞜����de�m�c���V��i�(�ދ��L�c~/�3�=`S����J�_�֨�-.��>���ۓ��J���(��EN����cou؇Pm��]�@C�1��7뢳�B�x��t������V��@�=�����yF�Ŏ~�[����������~�u��t7>&�$���A�3���|���$lH_yd�/Q'���Š?�H�8��쇙��W����I����H����� Lw�-A�`��Y������\I��D�$���3�=����D5��Ȇx���R/�[-�H�/�C��_��K�sy�E(�T�Io'���TeG�mn���.�� B'��9zE�G>rm�!u ^���+��&W��x���?�w�"8��2(��״�FԴ�,�RDŲ��N5t�״������u����I�d��XQ
C��r���X��
P{��mu�e��/��r�d#��O�	���!��B�j��BNz�{Iz�ֈGI![����w�G��,�x���ln7-��d��]{q���Zr�E��cnXw�v�������
����6_N̚�_����%��n�5e�nHT�-��m�)�(WX*����s�O�3�W��O���x�V���*ql}:|L�G�h��Yke#���}$��F��fg9m[����iyCm�� ��`]��By��r��,,&jg����q��).|�UXj4�/u�v�B"6<q�zr��u����q� a�u1b�� ���}�_u��}1qBb����kz|�UI���|��d��{�b���;�4�ԤP��,,b�����
�FC��f���؁olvH�\�~��l�J�x̈Z�3[�&�!��.�;d�!t��}-��1�ž��cJt	�˷���'h8�X���⤾�0��m�c���a���1��^��
��X.@�6�ߺ�I�p(�i;=P�� G���o���׸x|�-p@i�%Ş��1�k5Mb��Oc@�{$nt�OƦ���aŲ[p�=���EsY��G�����o�Q�`LL���A�����-ZM@X�F�� 9Ҵ8z�3!}�5f����Foyn#��&V�������c��o�xk��GY=K���C���;����oL<u�AP ��כ`�
^�a��YL��Х=�V��pvn{RM���^ۜA�b��#1����ͻ(����:�H�sJ�̸��m~@&��{�"�J�+7���{�����3�.a�w�V6��FOfi������0{wZ6�?=j!����5��^�?�8{�Ү!�]Y�e�,sQN@h�M�6?c<�2�1�ڿ�b)�|hc�\( ���k�j��¾W�C����#���%P��Y�4�-@v�'f�K�'�۠�w:��X���P��,0�A���_#�I�B�L�/�SX�;M�V�Qؑ�{R�lTD�(��YC� a���D1����P�,���  ��6�d���)�&	��&wZs#�W-7�&�*H�VR^��D�fE���	��G��:��;�v��y]��L�)�����*��n* �n�:ـw�t�E�S��Q�w�U������R��%�azy�x[�F�}=�[)��0�:�?K9�SQ_�ϙq�Y�gj�� ��v�M���-\�� &w�J�[{YoZžo5eL$�7:T
������/v8��@�.0>�n	��Wc�i\l�w�ZY.��Uc��L�eL�"n��TGd�jòP��~��Y`t���߆nx���h���*?i/���j�Ě%i�1a|� =��8j8�.]��P�T>Rӥj7+h�ih嚗��
D(Aa�7��un@ӯ�L�hu캒���ָ�W�G�8G�O]�A���\R�C̖S�FH��32�1$k�X�,ר.���&�d�1i�W)�(���.�P�����(}��A}�8؂��1!�g�������{�4ѽi,r� r���W��EP�$mh��i�YP6��lt�KC�J���'�@\��}����H�0jE��Ƚ�9ss�A���qP޲ĩw���ݟ�6:6=9虋������{�����ىì^�cU'S{#��4*��(��$���w�ܻ�o����m�I�ҕ��:��J�����r�B~#�FT�sJ���8jn����;{���I�M�h�-�a>��3)��\a&g}��u����~d�i�%�L�rԃXZ0}&�m�����u���](t@���=̴�������=��;�s��&>�-l��4Z{�����_�' fb�h����;n�tL/� Z��o˟��X<r�F-��c�%�5���N�Z�=���B�m�!�v�̼��I�ڡ�R
�:�9�}

�Յ��VM6�G�ڌ��H�.r;ɩ�8��O��]m�X��9ώ�a�Ͻ�0�y6.I�����������T8�$+$�__��@G$,C�i֟������nLki;�T	�%%+��(LS����`�K�[*���:L���s.����eJqtN'^�NQ���g��9���!J`��\�@/���f�#)�˰�vB�Q'Bܟ��U��%�Q-��"����4�-������4����A�����5���ɽr�9�A�����sJ�M'O�q]ú��)���z��u��8�}���'��Ђ���'��u �A;�}p�� �N�?�vE�E ��[�<Pɚ�:h�)GE��4��;o�# �,��-T�&'��d{~y��RRd����	d���]>8`˘^��o�D�F�jt�8��F��́� ��SBI��<:��>P�E�	#���-9����ytEh�<���T���d!
�9�}���Rn�Zq� 4�uF�.�+����}R�f��i@F��y���ˈ�c_�Dr��E]�zv"���&��
po��݋4�o���g���8`v�|�F�4����	"Ck�,�H�M��`n�8Ej�|K�\=�N=�<��!o�����f�S�> ����6�I��9Ϝ��=��ڇ�"�s���D�j%�\��:���r���iK)�)��ݚ�ƗQ`z��5p�0�l� �.�!������v�:�v*ؒr�j&�j��=}l�2׃�M�2�(@ãm�d�X�q|%��щ��+�'I�C.��J��q�CꄤQ6!w�_�'�O@{o\�����&��'���D�5�×L��yq�*f�5�L@c���=gk�nc�k�/ص�8w��5������ �N�P�N<2���x������ �[c)�hw�;LZ�����k��#�+U :�Q~m�"�,冝 ��zC�x0��N��x�����4����s��.��YYLz�����8�6��w��B�uzma�A�kF�g#g[;Ai޿��<u�ȶ���5ɭ��Ó��]��ϲr`S�3��JL�'��`��4��Y�OJ��6!?��
���bN���y���zV���5R[���w�= a���*����#ѫ�W��RV��T��`�I����QM|7!�]������`�;0�۷����m���k�􏹼	��qY9�qK��Z��.I����bȼ�Υ,�d��4��b�{%̥�Z��5���7�ډ�eHB��f�a�nT��cf[jӬ�~2\�����umF����b�e��Rd�64��y`݌����L'!k��J�h���[��������7yM�+���-f9-̕]W3���z_<�5�I���������#��͂�|CJ���t?�J?/������!t��jE'1�a��t7�)��]�e�(�޻"w�d*N0�5�O�
�Nc�h�6G9����\Ih)5&�"B`.��%��8a�ۊ5F����ji@��SCBN��Y�F���	���EV!�|���$��� �lSs�x2~��^T�;�pw�Pg��}~�M06c�^]B�o�L�P�I
90_S��r�������!AbE�S{�aN����'R��vbz��No|*	yx��Q6M+���<��G���`N����`�W����pU��XfaJ�.��w���4��k�l����yT�_f=��3�r�:Y��?�8�*�"[�y���B�NOK&��>��"v�5x+�3��ī��&�נr!h��,���Jd[��Z+'U]��R͖����� ����h�&Kz�}���ճy*����_?)r,h�i�/�N��lY�b��܈Q�TL��X=ٶ�Œ�վ�����&LE"�BD+ _��sMW����IC *Q�Hw	V�e�`bum��T	�D�M����;[�^xn˞']ȕ�qȝP�=>�Ji�qwn�!.�q?f�z\�C+�����[H}�4m���G�ry�c;�I�0<`�x]�)ɒY�5'u}�p�8��r3�џi�עgtޞC��5�"�?���Cه�,d&�<�\VK��PD��E�����!xz��{IF��M��b�c_RR�$��Ԭ�<�3.�a� �Tcv�k,�p�7���H�Ysc�-A�â�l��e���/���	;�?X�T�J�7��PE�Zx�W[E�曃=�MJ����Uz+�ٝD���P�[x2\�#�C���qB��}���.��<����R�L��W�����jb�hD*�w9�9>Z��C���>p�����6�����	��>4�C�bcR�h#:���/}� �\r?��5�z+�[�G�:p*�'�G<5g�Y�2Wǅ�ֽcW	������Lҗ_c�����l��%>j׾r@�/�/`K���n�+��r�B��')c�̴ηP���-����K,lTU����F�Z�Gˁ!�2�����9WؓC�q�����B���r��"�y^?���]��g/�$���w�&'�.�&�[t��&`�SK
��[ё	Ck.Q?�q��>��ft�����'�90���X�8�j�s�b�<R�
�[2/��#Ŧ��y��u}��nȒ*}DT�E�;A�����d�]��).��鹤�R�7��āU�::���`��:�)}#,�r���V�#Ax�IB>�/���e�3��[��6rK�ρg�8K7q��om���;������N T3�����D�`��V��֙����́�?vRdw�|%}9Yt{WQnםP����Bi��݉�k��)���M6�wQ��E�T��b��(��
�\H~�aVrZ-�k�t�>�,u*r\�M`���
y8eN��<��ŘFWI����a�PVX�Y�f��5,�zVYj�����@��-�fw���N���KmT4@\V^鱆��Z���%~��v*�u�a���+���{o���Ǝ�;�.�c-�|��?�5��8�d_��J�F �ۈ<%Jn�lI�8��Q"%�4�����䐽t� QSv�|���zJ��L�J`������
��Y�SH�w���yd=�7��Í�8�p�Z������C�'M��ǋY�$��nd�@juf-;���}�SPD�&�h-��x4�n��1�|H�jA��qw�x(0�w�'*Ò�1�ZX!�*z�7����t������[n]�H���݈��iC����뇉k<��H����ؿ�����-��4�a��=m)����͆��+,m������F��-8o����'���D#��:��S%*���kb�"�[\��¶����=�T��\��_��$idQ)+�����|���&?a1���[�rN�#C(�����슘�(V�n/��u�Tֺ���d�޶�BD�F�ָ�zT:����-��B�7F41�˙5ʜ�����/�u�9T�o�υ�rv�H=A�-��\ᑠ o"Bls��n|���8!�̀���E�m~�}�cDt����:���I��Y�����o�U��F�,:��a� ���(�R�Ne��*�"o�6�!��[�r��Wr��3����{�롡�8��t����	�g�X�	�F�y��C	��s���]�f��q��om��/�\�|F��^D�0$�V��%a�L��4����;ѐ�rU�3[���nZH|��"�����p�"�9��2�O��}���,~5�\o���nw�K��J1���P*�o��+�C�q�R�8K�,��[��0��2j�2��dL}��q�n%�e4�ǰR������@��lC���is�o��Ş#�:���YnH�����`��"�h󙽭�%A/�(��d��9��x)k$u�y��Q�t]����⓶��hB�����Em`߀�`���,N�/,�tU缩�i<���Yc#	h��sT)� *��#�Y��������b��-ԕdc�N+FU���������FǴeYf���Y��W�"l�HŹn䩖�
ue"#h��?�x��tQnk�Ĺp��A�����]����v�!��t)'��)q��\(N��d�����I.���^S���p�<�R_��x�b���ֲgC��&��s���V�'�i�u�E������Q:y�Ӓ���>��(�nz5nyK�>t���E�H��(h��&���*���KL|\�;��?�a*õ��"�D��@���q�{"�_����c<��:2@^�!f���}��/s�v����>�a����CH\.�.��3d_-Cɣ�2�('��4���ޯ� �aB9�H�9��bdE+d�k���?�	���ŕ�.�0>⬿r<�i�y��c�TcuA+�WLo�/��~�h�
�\G6���mF���k#_%���5V6�o >H��h/��e����-��)�m%S,cӞO��u2/#������wyo��c^�PM�L]��y��&঎%؈n���<t\B�8\@
+۞0�.���7<n F�;��y��7eD)�y�������¼�v���,Y��?��p�Y%o��c�����=�Td1�x�W�Bw�pTA �¿`�rz��TA,�'/�����9Bs-��]�#�������H�"��ޟ�j*O? ˡ������U�Z���掛"˄�'�d�v�a|��Z���%��]U����t��qݲ�˗ '�*��9u�����_=��l6D�ns����OQ�3'����.M�XZ'��v�.��[I3�H���y�ET1wl�]�������#��h�����p��Pd��n�l*=��級���lV��?�b;։�P�0 z X ��IN�b|�r��厀W�,@OD߾ڛ��?��خL?$1��x�Y:�d��{ڇ-��D����#FR�Pޤ��Og����]G���� 9��֌A�Q�ԍ�VD&���6��N�1i�C<�̌�i���eg(�n��*�|vf�H>B�T��bGu�a��0d92��	6�rp�N��:oUGr&j�Ǐ	gv�;�u*��iR�U��p��xo�V�]�Hk��}@"��~8`0GX]�����v�	g����x���3lF\BAd��h5|����#���Ə�hݲ��Ĝ@�-
3g�nW��"Ѓ����H:.�l.�W#���eO��T�SO���~�0�wX���������~{2��J�rAG��X�p��pV,��=\"���>Ќ}�N@dM���Kߨ�]��}Lb$�����댃�lΖis�&�摥6�7׎.�.�(ր�n��S�{|p���	�t|kϋ8�:�}@��8ϼ�;��x-;�_+2�it��.Oׄra��{�"U�؜F�֣�ІM�,E�l!O������ձ�F�a����\Y��8���@\�Z�ϔܗe�ܪL�[�����S�R�ܪ���y�pUt׮�Tܿ(�v��}|�����G�}T��qirו
�c�����'�
D��SB� �����Yl���|P�,{����ސ�-�g䋇�><(&�?��e��o;R���ωs��M�V����=%����w9f�KyrxP�|�o�岎7�b^���KYD� =���1�'����1�:U�zt���
�=�$�`�伨����=�0�ã�mk���z1�c�#�"��h�g�#�i��������̥��%za<��UWl����.C,�B���i2϶1�B��LT=Y��o�I�T���[ĸ�q��n�;Kwv��<7P��
`�nk0C7+P9�gw*G�6YR��r�a?~����i=R?�����
�fT��@�u(��,%9�n����|>�^�Pǫ����|���T�|c��&nI7sMr��2Ej��I^��+���a�;��A?��샛_9�zյ8������s\(4oѲh�s��,̄PO;Y����$�y_S�~W�%�Cm�D0��Q��� �]�.�][%-��CTF�^������:z΋�gw�A�JA��0��7���"�@`2:ۺ��§���xN���-�΃�Q�K)@ѹ��Ժ�I4\*�:�^��J�U��� ����É۳�Z�@�K���%�$<;��B�Lw?��Ρ�%V�!��:m�O˘�����,˘��~O�=���L��¸&_v]R�K�OC���%Q�������q�����|���0�
\N�`����G�'�D��/tut�-H�g��������B���ae�U@o=p����L'�#Lr�!V�u,���R�QMn�'����IZ���[���LLO���f�+��k�*7^��y�I+���`�}��T~�}q�)�?1��Z&斱�L!얼Л�&)˗�q����� ��b7��J����2�"������� Y���㧌�k0邫�h���S"!�.���a_Go�#�8Xb	�7F�t��U��x����t��p��#��;�Q��m�>U޽�ɭ�� SE���*xk����*�0�����褒"�:P��a�!�Ę���#|�����?*(���$-�0�ws�/���΃������9%�-8S���t��� ��嘕ݿH �	�z�16cPt 
�,�Sש���;.=�Y��P�墬-��~���<�1l�dl�a=a�`��J:��֧0L��T=�W�a��G��NI��^,�/W��Ȅ���6�kP�x�
P�n���A����͙�Ҹ��C@8�h�Wa���iJ�_Z�+����w֔�q֧:UÔI�Җ\�wHE�<2�x��V�fHjov��8�n�����1�l�iCܲ��
�=G�K<�����n2E�ט�!��uoEa�Q:F��N1{K�����O��q۪\8�*��8�{�B�f�Qg)z�;f�SD!g=���J\�l��A-�U��_���$�������X�7���Գ�(�e�NS����z�- ���A&��H��v�?Ŧ����M*ߑ�1��:T *,�鸀l��j�޷�7/������4	��j���5��[��kq�GR!���Z�J�s <(2 2��Ox%�3�t���K]Kh��d%t�|-pyl�A�U9�_e��epP�B�J���	e��������JK��z����;oq~	���XY��z�9��'_uA���N����7r2H���M��|'7���JA��2�Z�`���d�{G�椴	�߂�|"i�W���+�!��Ʒ<�����B��~�.�5�.n%n�%ϭѼ����kK�B��U>�An�Pkt�2�:�F���@��/8v\��kv�[�H����U,���;��
��^���S�o���t�b=4�b=6cS$���V���Hä
�|� X��{�;7.;B�+(�1M��{�°DC[(�*#J���!%r�u��]0�TJ��Z,h�{��;Z��ғ(,�#H��.= Y�79LR�:H5����3f?��[SD��up"��j�q¬���O�G,�e��J�҄gP��ӡ]��
�`�D#�
�ϐ��V�Bծw�<�b=8���J���Y�x�F�\\���m�E�Z�Ybh����7�zr�r�+6GA��s���\��Cŕ��o���q��5��P&��zw��;Z1]0����XM��0>�J�&?���G���ؚ�W{�~즘��?R�?��!� ��"ɀ���yVK�;��r��ix��c �I�%�cϘ�Ɠ��2�?ws��k���þ�S�Z5cH�Z���U@�V�?+Y��`��p\9Ɵ�nT)����8A�8}��R�����y�+�+\�}�{�ߙhĥD�A?=�$x,��:�;���]�-�.���9e`>�]%!���J�a�߯v3'u���H&����3Dհ��y��FlT#��p�5�H��=��������������#~�@:�?P��_�cpIA���)�3�MUXO��Jk����}��2�P�'[��N�������v�=��5�*�G���k� B���x�J�v�|#��eU%Uo�b!		��|^��m�odf��1�%*����~�F��V�����p1�*����Ÿ�/Aɬh�W�4�°�H!;��hب�9����Q��kQ�=q!�7�HQ���	�K.�l�嘯�Z�=��@����og�{�d;v8�6+.��*]X9��弯s�J}��^����W����^�v�NrҮ�3�'T�2�B�"`��N�qk!���!��f�|��m����o�`�+	���I�UA`��A�gE2*��,f�T�0 ~����[Z��ڷလ_�Oo3���~�RбYV��C�H�)#S���x^�}GZښ��¾aǄ�(�x��§H�{���9�D���R\-}Q���yiR�h�2!J�	~u�n~{��Y�P Y����r0u
(=4Q
"A9�WĘ�Ҧ锚���Y4����THv	��%k�b�~�ۼ�H�p�w�	r�_�6���4|5P���>��6���ۈ��<�&US��W�6�=�w`�|�Q��c�m�n\L�� �xa����b���5�>�r�8�QJ�>�ہ`s觮���OTD�Ǵs-2����O�.G���n��@ȵ�tƸ��͏B��f�����Т�I����6nf���̣4�JC���$��e����g���s9���E�YY�S[��Q-�Z����97�y�%��z��hֈ�,*�O�q�Ʀ�{|_m�SV̠ :�/�g�Q>%JhE|~�[���&�6F��A3�o4�V�8�YF]H,�0�3~�ezPoI�����Zk<k�ty4/o�'L`�-�C�G� �+gC�h�R���U��FE�0�5�H	�wEi��
u(��h׻����K{���}�_O.T���� ŷ�;̭J%2բc
�,�
��aB�T���G"nۘ�L	VG��yIx!\�5�ة1�
ev�н�agm���@��8�R�_��Xv� Ɍe:Lb��u������ʭ��5F����!�,�]7�2<u��%h厽y�@��c���L��v�_ͿSE��)3��䉲Հ��+#�,?�M7h_:9?�詉7��"�:��3��A�f+byR%�->TM$>K4��z/�Q5ۢl� ]���#S�ш�����E '�P�P#��і�R����4_�>��?L2^�pVg�U�~5Ʃ!���1�(�ǈ�S%�r�MY���M{�\��Zɰy���+"�ցѺ<�V;���$U�#����J���V�}* �@O�~\8��1���'hz5�M%ue�(Ttf1$Xm�V[�G���NX��b�d�hN�]o%3�@�>
<{[��m[�Lj'wp�8p�݋��V��MM���_҄JEĦ(�d ���ĉ�VE.��dL-��0�^������uc� Sہ_Y�bX���ؿ���l�p���6JXnq�[��Wk�=#P�$�ܛ�ǁ�_�H�����+!��d�:6V��/��Vw�`܈!Բ���K�U�(�3�ÿ|M�3�a �l��N�Q�����.S6��oʉ���X���D1��5�ő��a�4��࢔U�q��W�ԓ#�0���3
r�h�ܔS� /�<���8^�5#_l��FS�B��9NS۪���m�0m�ъL�.ڶ�9-jߖ/�ǹMu�VzR;������j���y��Ɛ���������_�S6��)x�y�)��V�~��̢aO�þ�}�cө�|������\�Ia#����Ƞ��L>�h�:!:��F��j��A����1���ER6J䞔	��V�L8�#s�P'��2��`l/"��k��,W ���n�}~�%�mÏ9F!�����͊���ԃ�Wj��G�)�98�͙D��,�x6��%=�!0���~��J5&G��-�K�PJ$vk�LPfE%�a7�p;��kKDy�dE�7���Ss,Q�濋/�i��I����/�,D!��t/�(0Cl��MБ�GZ��J8U�}����o����ֶ��$9t��7�+�H�Wń����
�|��%�c�k�MF��*@Čg��6�l����R{~��'��
b�F���׵y0X�L��> V9�����Zt�i�M�1���.W9��DB},*$����o,�����E=�iդj��:%�抙�#h���-�����T�]�X>a7��:b�^'���WhZI�}�CC����ꥈ$NVi�+��^1���4�bF�����=^ӻ*V�����<�MD�m#�A��~%�L��U��!�l_�ӓs}��1�3�l�qj�;��f������h�!�����R(c�k����2c|H\<��������F"veY�R���?[��������.�St${b�BS��et!4�b�����n(��Џğ)��'�>`��ǃ	�(Y��-m�G�:�Q��8a�J0���-%g�������EdC%��n��+�ʊ���e��-6��X�S+�����+c�i�.��������9�����B�(��V/�s��*��i�	��<ݰ�.`9�	�W�H:Azq%��!|j��?V��H?��4:�X�xw��3�a��ڱ����,�������㽻���vg׈��Y����S��7�=��v��dC\��~�	�YyQ����<����R;a�g
DVfV�e��HIi7�5�dj�8w�	9�� eHh��pq��+YZ]��{P�LD:*}Yn�v?�:�U�*�KU��Yj��)����g�=�)}���v�ӎ�*���_T�����.��!p�z��聝6�P���l���g�y9���lEPn1���5�%0q����R���YX�_
��٘����@�~�VU8�~ ��9��G'�K��+��P8�M�wr'�^?� rc����G�N���M������\�D|ä�.�L�����y��z�w?��+@gS �����o>b�Z��dm ��)7�>:�Lj�:����-�kPb饊F�k I`0��o�nO�B�\�Ü�0��s�@q��^�6�A��tV�>X�*�#\�;w�E<��Cץք�ѭ	:Ҧ�~]W�G��*���&Xwyu�N����&\�=ߺ���&�X�7��ʜ�lX�榁��1ѣ;��ȂR�f1K���k� ��א*L���p�4ӣ07H^,�}W~&��.EװԩWB�g��z�0q/ �T���3D�
(nF��q4Z��"	M�K�uW�n�79�D)D�q�*�X�9|E�,��j���1��P}�ͽ���,�rq_`gL�>t��L�y�������itҵ���ěM-�p��K��AB�Wr��O�&�,@
U�uaK��\k�z�O�;�I�Lm�F�ZP�?W_�� �^�K�R���l����cD�D5�96��R�K$�R�v&dӲ���e�"!Dx��I�_��g� eѻ\��G��^a{����t7[�� V����,5��~�/h���R�������<���A=RQ��4R�a�[@�O�`@Ept�`�s@��m�p��@�19Lm׋���W���ӌ8����\=I2���Dk$La�W���ỷ�]q(k|4����ؼ�U�\ ��94�Q����3��;OFN{Lb.ӏsN<6�f��[��*t�
b9�O�FV���q����~�\9�v�T}W��W��8	'�*`��2�������OB�C�̘����&����J�E �R�YE�%EA(�%#$�Cs~?!ny)�.��9��g�/��E7�yg�a}�ʕ�s�4�E�R�Q_܃�p����sl�T��݋5���ѻn[k�Э���I��mR���.���/n���UȬr��k�����(����R�SV�^v�p����(���i�՞cN�F��'�7����-�s�®G�y�D	���_����f��Q>ʔ���^r?dd��B�W\̛���1��5��)�f�O;/�`ڛ��q��Z~�(k"��,�s�@H:=�\����
m���M܎��ޗk7ָ�R�(�K�?��*��\f��٧CX�4ˡ~�q�8��M�Jv�G4Ar[W���ȭ�m��S���>V:F�]-M7�v���RzP�;�ȺPMW0��>�ŕd�z:,�&"��4 C]��En���o���W��)��$3�XX��=��/3��Ų��z��e��{��q@3]e僋�_8E��s�'*�/��i�����#�����2K��疛�1��CsE�5O��D���(�`������=�#�懔X(r���p!���V���o�몿�>f�`�`U�`#���.E��2���j(�o�-�"ׅ�b̦B"R���	���?>����w�m��C������:��&'�<�!f^�T�@\j�	\�H&/�4Ԑ?��̾x�\,�h(b���he�y�!���]8u��m��l�t�\W�\R;a�gݎ�q20�6�!G�"��פKs�r���;q+�=�·7����f®�<���J�b]�D%3���,r[�v ���#���KY�����	�����g��}I�[�VRT?.�f��	�Qɻ���Q����A=�3AZ�	�ʏ3лeW�X�s$��Ѵ�f�b,s@�������"U������������%L\˭'%�\�l[P�ZS���V�+�u�&:#���L�m�D=��mUw����h�v��,b�j  5���-U�!C1*�"��\�����1r.�re�������K�z��rz�I�Ӆ��N�i������n�����&�Q�X�)�|EU��ҹ�%�������$�����+���?�u�Y��Ɩ�̓��G�ڪ$�	Ue���)�+2,�n�@!a�_�ĝ"�7��
JT��O;\y�X�~���A��L%� ��}!��ܺz2�3�"����H��>��l`��a��Q�-��FDwG��kkN7T;ٻ�3;��F����р���ǹHw�Z�A����E��Q���)H|� �W���B�3Ky0��\I�z��/a#yE\{���Z�V}��j]�Z�4I��75�X�Z��3��j��4
�C��e"qז� pJ��o����L���]+�"��0f/;Hy��1z��w��*dY������B)Ǽ#��߽��{%s�K��1V^�	���p����S������`��Ǉ1�L�/Tj[-%��Ϯ.��-��)Y\�nm��{΢�.��1Kz��CI��3��y�%(��^�P�	WVU�G��+��=����<��Û��� �Ѓ3͟��z�c�;K��,x�4a�ѽm���h��N��7f;+2�%!h�o5��{��vT��=�	��6e�-�X�������ɥo�B����@���)�?��%ƥ.3�(��S�t������c��	��������e%IRD0ïxȔ��h��A6A�W��F�p�h�����������{�ke�����T���3?W�j��B��R������B�3Z��By���h$8�?s�Bmy������"�����B�ٞES�����6ʜ������x�����7pa��̥�>�\@a��A���(�*�#e&h�0��6Jr��i�`
O�[�!��LZ��>��P����@8��=b���{
_�0;M˺*䪰z���A��X������$��v)XP��6qI<D���mp/�������/���	D[�Q�i�bu�((2ڍ
f��^v2�Zy�-HN�C��	��~�<B&���q����8e�k�]�.g��ڲ%󖕫CK`�l�#v��l��Ʉx_!�����H��쟝ǵ.>ǥD��h�˫��*��-��A�C��G8�u��i)��@]���X���C��!IE|T@���a��V
��M1���(zM�-*G�>,��rr�ھ��R�h��R_S�`\?*�%R}�}$�/W���w�l����+�G L,	Tp�c)� �{� �>�pZn����D|k�ho�Ma_���f���A'%�0V�FEw��3I>4g�]�w�sp����q�߽�W����3c��A�������ȶ�܇|s�*�6gg�I��cM�Gk�����O��j��J�����p�ǧ/oR �5��`�DOl�k����lPa�:��F-���Tp��m�Q���U��=���Tҋ_�齡���w1�R����
�T�*8�V� O!�_���bϻ�T��{+%�Ι��#��9�-#-d�<�蔨�A���x�͖����8�ehZ��x��i���ܠ�Z[�6+7��0� z#�
�4�l��v��U�ﭫ�d�ƫ�Ԡ��N��mw7Ӌk��l��;�-?\�!�zR�.5� ��Ȱ��(�z���x�!��N%(�����h� 8����$��m��u����{�M�[	�F&�r�=Q���bY�����S
&o�P$��(,r�%�~���Tx�0�t�6��D��Eli�.܆��ī�hmi�O�LI�U2����_L��G�d1s'!8�~�H������Тf_k��V����o��y�7������*[��`;�u�6���V5���F=[粖,/�8a��Mz�嵀(qn�*�L���kɜ�c���[���h�~A_I����P�`|h�p��xEg�׫?�0�Uٙ���r��TA�kS�oA�G�)��ή,*Zfʏe⑰Å>iOgޒ�v���o���:_�0ũE��J�xʼ�p�����u�`����x΃��R%����b̓�yg'.�au����%#Ca���j,�uX\Ns�*;|v������x8Tݘ&d�����2��� ˢ�ynɵ�S܄GF]��V+Q���J~�J��\���]��X���Ji����C�,�������ؽ��S��e��7���E�������|�!���s�"�7�H�/�$�([X��0��׈�������ɧB�͹Y�Q3�#�cZ�E6�(�DTnZrht�pP�&�7ڭU�@�&T��@� t�Ƅ�3�N�ɗ�3�2�������6!���P.����-,���|�<�D�E���9JjN �/^'!�r�hq�ޣ=p�
6=V���G�&����Y��}GH5���@A��,B��e8b/��O8 Eh�ь`�.V��������	��G[O�n�]��
��6���,�ʟݝ��/��C	�!I�+��t�6�]�o�B����J�[����_�S���c��Xm �KI�����m<Zd$8�� ��lA�n��yS��ɿ�;y:�`P��?7v?Ş�ssb�a\�w��q�#t\6�3����%�@�u���5Y #	�z�ػD���F��Y|�Qj��m~߈��6�m�]^�/iV��*�+)�R=��5���L^����]I�cQ"|n����+���5��gY����������u��M#���~�s�Ѵ�j�t���w� H.T����I͵��v��R)=�-��v�h�gO�����2־.��@�/v7�FS
?	qQV�F�Y��: �W��|�'�s��d�z�k.����*�, ��I ϰ,��mýXvd��ɐY��f�� �
��
���x��I�c���31�h�M�'���u�4i��q�C�[��W�_c��:	�67J����+x^��>
��-]. ��Q|�Y��t]f�`sc�axw蔪�BJ-�MU����*���$(S��c�\�>QE���	J�8��J��F��˰�N'P�a��瓸IQZ|�� A$����|o�gW����o�]Ncwr֌�!�RvW]�aM�A˖��ȩ�V���UP�^>�fK��BKXyRL6C��^���l'��,¾��)��hO>Kv9���
��zU�H��k��*���#;��UtH�&Q����<[��J��J��|d��~�kպ��#�q��/���+9ïS�e��'d���"�K����ɝ�+D��J�![�㒋���-����(!��v��@}EsU�v���jy��p��=A8���c���3�ճ2a�Eb��`;n���@��j:v�&���B�GJ���,����w]$��o��Q�����eï�!����%M�����?:ι道�[n��w���=�lH����a$I��V��� ;�V�Z��aK�6�|89���(x��HS"����^^%�H�
2�?a/⟯��ꃎ�i��\(��#>�pc6%��`��	0���RP �F�R�\<�d�y�Z�V����D� ;�zz	�Y��
 �$|����u3�o��*�Hz�G��,|��7}��D7d]���"�L���j��&Z�J*���x{]}���'p�F�E䎪Jd�R�L;[�F�C��q>e>
���܊EzTO2 %�r�m�﹝IK�2�*I<~�cEd��dg�0Ok �����f�_�J&���g.W1�!	����dtw^�\� 8a�~N&�tJp
�Q�)���$�c
1ﴀ���a�g�C�������߱8�����T���S�;R�j�$��8a �|�����?Qq�����8���h��wx��T���:���}!���~m#(!�Jj_"n�u�k6<���F6D]\C�����	�P�G�
��B}m�)�^�0M�\���L�=�$�}�E�߼��.�oVt�lw���@��z=������K�:���z3g�jEB����<Ya���=L�!�{��̐�'�c�y�S~S�����c@/拿6��>�����lp�Ɠ��P�4���QG��`��ߝ��a���0���8Z'��Y����m=�.t��nU��z F�����vE|�~����gș-�n�k�&9��{�>y4�qm���(�L7���i�l�'aj����zt�Z�3��
�Z�v[��3��-�>��6�˞�5R^}7�Bf�%�r.;*X���"s�=^�;�uk�"�v��7��-k.�$6.6��Ӧ�K�G����g�W&���9bL��r�)�_��_ ,�ژ��M�T!#���b��{����"������1�U��'󚱑���{�W��n:߬����q��|�v-�z��V���P��X�V�D&yFe!C��ٙ�N{�]�S��9�]����b�dc�;Y��-�8+չZ�G2>@a��������,��`�g�~t	G|J�C舘@FK
���M���﫳>���Y����b����b������ȵ?�Bj#�o��J�q!�ы���{�F�o`k6�{++�z�Z~.�W����g��*a�z�Ț\ܗϥ劝W���f������e��kXX������t�x�!�@�g~چH�~�40[5'���՛�h�]����_D9�q�o�<�)�'87xo�k��� 明-�����r�;��ސ�Y9�7;�����9�܀H��Y@�H*jc�D&~�UL���o״t��&�{ud��:�y #�A;�)V�B���k�r-f��H�gZ�C��8���*�I�_u0�כֿ�zҏ����K1hT;����}4����*���Dқ��h_��ptt;�̳���F'ʰ�[4����.B6d/��w��h���f�ۊZ���?�2���0��2P}��&koJ�^y��,�
���Dm�k�Gz��~�A>n�}��y�d7sޫ�b�VM�}�`��S��t�t��J��S�7N�꿁ⓥ|kȯ�gʘ�-����������+��G	�(ڒ��A��h�G%���n��;�1��ZT{�<�9l�	�>"�}�d��;/c�%��a8뾋�G!��;:��� l��-v��g��>;�[A��3��TK��p�%���&<E�@[Ә�I���e%�V]v���	���UO�*F���p�J|���{�Nlð�|y��U���x��)
��0�����:�����w<n�e�+ɸ����
f��Yk�<�dub�#%zz�n"�J���y��J��ӥ�[����^����������ՙ��/7�y����R(����O[�i' 9�e��
�)���_p��bF������S����9���(�>�����`�dzQ�1/�{b+�/zf	�FĦ����2�
EE�ǚL���Z��H��~$h%��۷��˝�d��V�����fc�I��8�gAr[���]�
6��ת�C;��[ohR� u �>&�D7����?y���od=�s��K�r�5߂v�
���5�z#L:+��$�5���rJ�]j������D!m|�>7V���ZEͬ�].`ʼ�����R�OE�l��6!	]姩�r��a��|A��ŬmR0��g��8@�œMD4�k^bU��9����K��/�	͸��_�o�(2aa'����������ƑVs��.5��2!r��'��4o+��֟����*�����OY�sͬ
�
�A�z��oģ�D,z�"7]3�
��$Y��_@���بD�{VMD���x���Q�����hti��f���0�@,���1��s�9eC��8���+Ǆ�0|��e�������yd��+���X����z��-[ɜNܟ�����U�m�M�gy�y��6S>m�bA.���ѭ����;g��	7y\�~*ʯ�SK �S� ������*l0�E���O�ľ���m��-� �*+�{�l�|j+-����:�)-E. ��7��B���
ަ�������� WƑ)aN�1��R����7(�0��n������?�ѯ%ڰ����Dj��2�zf%�@s��N'����D6�<Nj��"��3�9v��1��@�c�&��0/嘧p?R����G��ʽd�`��������Z+yтMoڜ���;�C��$q�lk��#~06�X���ړ��XW�R�U@9J!��.ZA?r�z]��ˠP߻��2�Kψu|�1��M�徝�w?�D��x�#|�~�;
t�XQ-�iA���v'������B�>��������N��}��{� ��H y@�7ȷR���x)��ρ���:�b�٨� �E�ɤ@v��#9���J92T��Syn���rV�8�d������B���!'�]JV�X-���B\f�n���^kƢ�=x�����V$C��-%��M��H� ���*�#<��q��*fϬN����#�v�,���x/�9�pz;;@�S$��o�a��w���?��ӭlj��q��řG퓺��4BIh9<�p�+�gU%h�b�|V�4TJ $�$�tL�;�;#:m�zr\P��c��u��S��BW[,�s��5C�E�mg�4��{����&�sW&_�����l��g�ҮgO��1^����,�rbN!���0e��f����\'j?������;T,j��A�����Z]�Z���>�*|ϨzװS����d)�Z{�oZi��i)��˦<٦��,�$Wγ��� rƇc�~h����7�|g5��8�-o �g��#�H�ϒ�����W�	���FS(:�!����g5�1��v,t�i�\��+�H%���7�z��!9��:���v\U�G)h.��EH��do�nn:E�Մ���Z��`�4)�ܒ�G*
3��X��&��J�x67,w-��q���ٮY���L�{�q`�(�:�t3��Ɓn�41�@!=���ک�BW�p�ytG �K�M63|�"8�Q��Z���+X�o��Q����7j�]ӡ[��a������3)-]Y"�� FZU�}!��똂Lp�ڝPE��;*�Pp�����Ί(�:��K@0��%�{@ufJI+���[�O���U�᪟�i󿊃��a���0cm�3�b up���n�6�_�;��Y�5!�H��B�mS���u��Qǀ�������@���{����\�?�F��"�O-i7q�d7�1��T8$�����1�MDWP�B4��W�j��f�"��� ,6�Z��h�T�Y���I���v���Gm_��序�9Z�v9����?3���Np���o��n�WǼ�$�чO J�pC-͟3㨤�����
�����x;���+��4j�����)&�9���p����-�a�F�p�fr����X��}�X�3D� ����[^��fAcpA-7�,���n;��|ODk�M��|^��ϑ�b'i/�W��?3�P�ߠ�� �^��M���j\���rG���g_b�_^9��eT3fn�<5Y&M��W�P��b?�&��NuX��HtN+�_N��/Ɛ� (*ط̇]5|�B������sy��aݏe��j�?,�i�.���>zH"ʏ��?>�bB�A�Jt����+ԭj�`��;��kΙJ��2��4+�����0 K�?�%��I�I�Gr99��>�n3�?q4�#Zc�/�+�l{��Y�z7|p������������E`ٵ6vf���L�&KӜ��H�6$0]� c��YM��W�'<����FG��b���0b���K�V�銢n� ��P�f)� >y�݅v�.w�}�˘�<��5*��|��� \e���_��Fi������~V
wp2�����i�M�b��9<2p,7,e�6��sr�[�t�B��k�&�p�Ag���@ή��U�^�:����
8������,�J�e�\�8B��C!��*s�J��h��<X�Yի��d�Fy��+�6��9��K�"�Us��K�g�
���ӎ�ڱfРs���\��1Z�[k`��*��Rǝ���I�i�� �1K]��������f����Yy�a�a�i52�e��T
y��K��6���q��[�Ӱ<��u�C!p}����@%%9(|t~�ȴ�{sv3�|�T��5jt�JΙ~tҿ~߼	=x��>BGʤ㟹���8�n��)�3�C��2��N��4X�dw?��}\B��3E��''����<a��Z�V�˶q:����v ���"`��ah-�`�(%�+1���[�T�u�~�����}
޴��3�pIu?�.��d)�֊�Wd&�,ϩ��>�W��%��'��	�Z�����~Ƣ}mE�T�y�eKR�(L�������	�y��������
�n���ҿJ_ŏ��@���'wŵ�״��j��#�(����/YA�- B�]#�
s�b3^0 [i����� x��P��=�+.�]e\�M���T�]��i�x:U��YA]�yJ� CY2�r�
V�(@�x{s�p���Z�']A������.X[ΧE���52%}���ͩ7��X�t��(U�;=�?��3!"�OH
�T�L�HJ����'��u;�+#�*js��>̮������4J��v7;�tx�.9.>�Q�[�`-%i1�m�F�D�ZcG�K����F~*�py��vi��G%AC��.��+>M���{Q���޷�R�e��k��1N�&K�3M����K���1Vx�Rw��ѐ����.��p*ۄ؟�r���jB�O��n��V����`�:�b�w�s�zZIuv���a;��\͡V��5�-�f�x�&�$���߻t+J�U�rc���'̱��ax�{��#F_�+��=zœ�����=�#TY���$P��/�PK��`N�+�I�y�zi#�b�GK/YKs�չ�4�Hv�4����|Ό)q4�z�+�oڥ�)�F�N�ʶ���F�'Œ��WC/X�E�%�>�ۡ�@��Y}ga��LH%��t��1!g*-�ב��H�j�
�t�}>��{�P4_Eb���.�GQ?�XT]%� �,�h�!�e^�'ov/���a�[����z����.K/L��5	�>)��W/���x�!�zq{y�i��}�*M1��I��{9����@�t.����'oG �#U��)j\<+���A�}�-f���'G�ƣ�76%`"+1�7r��ky��F�y	��b���I'{g�J�G���X$�̚�e�i����69Ƭ�S��IL����֣�����}�l�_��I��~���%7#���_�\�3��spL}�/�o�{7�N���{$�S��V�w������k�%MV/�n��J0�tљ�d�ͯ]�h���Dn���'�^��ʵSym�"�r�)��=?@ĉ�����l�'�?����v���@��x}KP�W�iy��D�Ao˄#�eLVm�N�&�c���%�A����vMр!g���v:�F�p�Y|A=��{:�^.�1�
�z��?�=�5{�Ƽ2��$�A��ʀMbмPUq(��WKo!�w+.d�-�2�-s��������:�B0݇��7���\������s����`��Q�� �yV�X�s� ���qNh� r�k͝7��l�.7bt��6޷u�-E������zX���F���gz.o���Lq��\�j��<�ۨ�ͯ��R�z��O�pY����@�_�Q�XX�s	�g���0a:}6z�')�N����M��8S��T,@�&7���r�i�?=�uY��Jp����e���W��P�M���Q73|_���JH�b���V�1y?�@�@����� 5�0��:���"�98#�.y�B(�}Յݬ�&F����н�Vg3r!�o�f��"��x���D��vHe�o�I�*35��$�`��)t����ܘ��44������S�������j�7A��W���O;Vb�
�:�8�Qv���Г<��K��q}Q���	�%�Κ��1��[�C�o%5��K�Ɉ�ZLklqB$�K��}�#��A����~i�ZV&�͹�bCd�����Hn�[���MJ������T%��(�6^ѹ瘖9��\��j�B��~��V��J�ԛ����|��Tˠ����. ����|4�Bm `� �mIQY>��Fn����]g�W\���F�'U};�Ӗ���n���!@�������Lr5�'ꆮ���=��c�ԅF�rS\� �͉Ɩ'pi�e��ۜ������J%�o��`AZY[��ǌ��&�'?h���IE(
��v=�mK��ٰp�4���EAa\�5�s�'G�đj�u T�A0�����٪�A{��OoEpT\�t�{���0��Y���e�4�pS���\i[T��.��V�n 8�eW�v��#QZ}�f�A �\�*�o򻓙��݊S��=zG�^T�1��H��4A>ߖH�� �����v�2�"6h	:X��6'DA�@@C@���Dd��~�D����V6�W�z�����=r����a�V�h���m�k=�I��H��6�B)�%G��O��͖�*ݴ\p��:6%%tB��ǰ��Zq�f��n������v�2�ƶ#[�e�ޞ�؃7�P���i ׀V@�șs��?��AcO��V��Tќ�k;�E�W�����&�N�G087�i��$f\Ę:XWk8��? ����(/���m��gᗡN���O���P^����K �_O���l����]�U�z�&����u�s�� ?&]����R�nƒ�M{a�
�Ծ[�E�/��/�t����遭�Yoh^�IZ�b�C2���� '��˹�	��
<u&���j鮡�I�F�a�t7}{�$z�"�rPs+�m�X�+�,�����A2��H6��^�ؙZk��f�J��No�`a�ź�:[*�h{	��r�񌯔�oɊ�m��	ƻ�4�r���@l�/�6�"��_��*������>�$��AX�Yn"<����r��#rƯ�nI�RJ��U�归�'�F�X��p�Kkz]>bm�iِ����a��>~H���mg1�<7ب�킋㮌8�↗��{E��q��v�2�
�l�4HeyGڤ�]�W�z�ʁUi뭄����u���:�fY�w���~?~��0;0���`�^��#�I��� ��<1�cS++���̡��Z6Y�8o�v{a�֚�Sr��`��p�݋G���d$IG�4cM������I!�4��K�?����"4��e�.IjA����.ze&�Ø���PJ��Gx���i~��i�>�=�g֮���e Ѫ���MbT�S ,G��/��Q���OWqq�!���.|L�/�'ѷ���|_����>��X�C�u~~5�x�.�}�JJ�ED�H٬\�%(5�eV/�GB��^m���c�0jMr�D�_�ay ߑ1�S�ި	�c�Q��c@��>%��C65k���t����
�u.Ҏ��魪>؋�W3|����W�g���^�N�XQN�3:�{uf'ܔ�	�����rW(���wT�O�W�D�xh�D|CG ��X�	̤�'Xa-j�`(
.�ims�A3p�a�K�Q[`�����p�Q�F>j
�lM���W��_���h7P�`�GR]SSm�U�v�9!��=���2e@O��f"�^����![ɽ�c}��'�� x��_EE� Cke��z"��o�(];K�����O���<b��DJ�x^i������
����j��b%wݨw�,���'L*D���4��d��j����l׌�Ȗ-g�܎��� ��Ij�&ݛ�5]ً`#��;)����|6��ꓬ�>1�̌�u�Q��ٮ@m^7��2�a�b7�A��̹*I��
�,���=Y�᭿�
i2���v���n���$٪�؈��L�.E���|x0���7�*M<}6���������J/QK%w}] {�=���цttɸ�5x�pZ2Gv0�6U�����8�������[�/�"��d�Y���(�Jt�"��3�y��p���g?���	�t99���]�4H�8�nze�0�u��7l��2��c�.�a@����i��@�Q$ *������nt>z���X�|�r����c%,�	��d��?��c=z�⯯�w����y�	���|�����YD��,��mO��_�8�b�K�pa��?2S{f�F2��^�n�3M]n��	<��X�C��s�!k 5�l�f̽�+)	רCY<�t�aF����[�ץ��z�Ғ�ZS��EQ��������~	��̐��_ii$5��n5@��Z6V'An��]�\�iecG�T�&�q�����E9uK ̷[�K���4Fb:bF�T��ۤ�U	���t�pEn'K��X>����m�(/3Lv��	��H�c�@k�mu�|����w�@�ez�p}ܒ�2_�3��qv<Q<Ɯ��b��K���:������*�G=��c�<Y��-��(*k�(�]����>Vr
V��i��=��+\�֜Z�8���c�j���%2�Y�`nW��ʑA:*P2�l�_��Ru�u��'��=��@1-ʞ�3��	Q�c5W�Tg�M�˸�28X'��R��t�q�Q=��^��S�S"��rQ�����H�I���N@������ݛo3�q�[ma�ݱ

�Z.~'f��>[#όwe�9�ʬ[�뉞�`�_Z�Y#�V�����2j�A��)Q�1(+T�'�+խq+F:W@���F�������T�`���ۮ�y���/���f�"�Vsµ�ȅ1�{�a�^��=�Tk_�{�1�a���c�2�7:D`6�5\Ϙ]R�6N=:�k>�,�ƣ�Ao/�4��-孻>�v]�U�������p����jq\?�V�(���&=��a�=.
]j�� �Ĉgto�S.W��mL"@��4�^�
Ղ3�B�j1ô��Y_�����C�T�V�0�1	h�IBT���/�
���W�4+�3e�v�N3��h�fzN�(�'$L��C�+7߽��lGfH���R��p�^�Fw�ᑖ8GH5M�倭?
ֈP|�W��"r�49]��j���w7�Ȱ�%Ρ(��;��k�7?ŧI���/`�����W��X{�E�J�e�?	�\�Ţ�(h؇0k��"��yL�rEme�H�g�U�_[	�*���gG&������;y��@�	x�*�)kD��	bH�R�;�z�>�q�5]��H�B���~�� YցA�*4�j�\�<]`-�OC[��2$�/Xk�|!�=�O��BA1�4��H�8U�&�/7:�&�UrM|��V�B�J�^Ğ�[%�e��#���E�x+���=im� ��a�1����+�8%�7��퇋$� �T���O;�i���R!�^���v�;�%� �W��s`�ֿ���K8Hf�D�B!P&��<ˀ� 
]u��yx�����Pb���`t�������o����|�o��S�+ǜJPje�	r�}(��S�3�:�@��a*�D"�LQ8����B�z��1�{����Q}��t�ӥ� �RR�X�O~]`2�s��<|���$��:IwNN��&�O���lnMw�޵�����G�i_o0���'XЬ7���wk��0{��I��?����Ycp����.�A Z�\��[���Ʀy�DƳ��D[j���v�� M�n�q����Ǵ8W?D�K�k�tlK���H�a�gH<���Bz����&-� ��	��w���#^����]n{��~^�8i>עm�Rʋ�hi���p���/&?�꽼����BaԜ�� ܳu��S��r�L'E{���S��J�ˆ�0�7��0���4�]G�R�F�7.�r3#�v���~!ݱ��>1z�^���T������^�1��dZ�A.߻O�7Aǧ�k�?�;���X,��=���|
s�ZC�i�x�\ �������|�XP"$=:Z�0ŊnE��
�2�o��V0�h�]-�8�Ȑ���e�S�F`�b�I�2�T%�q��_k�=[R�Y/�|6Au�Ho�S[��0J�AHDlZE/5����y�>��A�������$��a�d�N�����Oq�ym�`�q��'zrs/�'�ˎ��pPT�����?L�%��QDD���6Ah�z��(��/�ՠ��5Q:�R�-%	W��O�n:��H����]*��d�*�|� �8�+�+O��a���_c,&�Ge�iB��	D�H���-)B�_�ӝܲ�M���Z�џӈP/�X��YW*���8�8ǉѶ~��*��	.8�dܲ�'1��O(4W�3�����	�O���%/<��{����:�׹>~����v�!<f���7�{u��{'�jZ5��ݡ��릨>�F%&�>�IZ����1/���V]u��f�a@y\�����W8�-t�%���R�W��4��^�I���!:��5��7\!�
���\���6z��2R�v�y�g/#L��Z��?4��I�j��[5�Rc�𓺺��g�#���0�I���䎀WWrL�pN]�Q�E` ���d��7��"�Irr�l+�
	�~���)�)ȼ��Dp��>�g�~3�xD���G9s�O28A]ܧ�yO�#_��"��*���;�&�>YW���t�q�A2ߎ�ma')�:�>i�ȴ���Ϙ��a�XG�|V3�.'��}�_��{�����{��� d �D�,��-��\�,G竘�qO��?8�u����7��<g��!2�JgZ����w㶩@sn�#�O	#0�7��;-!*�������x�:�N��+u��G�Ž�)��҄��In;�*/g��F���WJ�w!�L�Q0'x�(��'xrH�Z*�8Ia���Q#(©�NX%�<��	h�B`2,�-�?ϛAbL�\���=0��$(����E�q�[70"hg�T� ��-����㊋/�GMD7�:1��w����P4�6� �5���UI��Q"y�,>�->��Lr'�O�T`Y�͔,8>���ek�m3��4�8�Y�6|v���d��h�ѓB�X3��nr�p�T7�CT�����ή��� 	iu��"W/#�^���\�w�>��6#2�N�%���f�D<�G���1؞7��)�ZS��:	\)���"��@�n=j]��SGm8h���i���1u�o�-��A�n{���}(��U��k E�J�� �AP���/�������)�]���9��T|��Zzk��Srҟ�.����)8l�ߴ(U(,q��Tk�j���HQ�R,xQ"f��g����*�
9<�7�4D �L��i�L��*-]5p�-H�����@�	:Pp���ot��_s�5���"d���!0<�l�q��R����1њ�d��D!���~|	�!w%��(��w[�M7��%zB�9=����=\<+��M}��o*�%q�d�+ή.��w�w!��qx���1��`پ|�e`��Y����l&oh�E���2��=���B�{���$�sO	�����_'��9V�U��S������6�w§��Ȑ��o�8�=�7](�F@�]�D��;��~��y��S�����*���U��T�ד���oC�~>��3 ���lr�R�@��M�!�8o��?��x�D���ėy/gw���/Q�CU��A tu�uG��/��/�V�(+���Ǌތ|���}�o�l��t 2D>3�!(�m̸S�������qd1��1k����>}�V\۵-?Fj� ���d���h���[�p�����z���ȋ�����ob8�h��r���x�1������#xj�"p4�������Dv䨉b2ϚJ�>B�͗���n�����~���y�}D�� g���GU�T�����}'s�B���-�z�1�Rf�$J�\�����{3�χ��Է2d��P̫��ˊ�t��;� �۟�W5�)�]��I�PJQ��C�(��������Xԣ�x.��9X��n��;8gY�N�'J�i��:�-J�~�,��8L8"@�ڔЃ̠�K���;�tP[%�Z/u��¿v���b�4$Z؞����b���W�����:I	�6��?[�T픞�Qţ��o��-sT_��yYʦ����� �7�$���� �zM�~h�X�$DU�8>)N����;u�x�슜���E�?�' ��fٿD�%dܷ�A����rfd5;��� Y2���h^�Vl���'f���@$'��
K)nr
.Ʒ�d��I�l!f��}�\yQ���[��0�)߳۲�p�U�A�a��"�l��T,���S���?/9I��sz����*���^�(�ɼMV��Tk��hO���Lɰ�C�g�V���_������ܿ��chZ�����;��D������]�Gz�A�n�[fx����,5�ձ�@��K�}�@b���b��D2�����p�m�[@Q���ĀgÁEF�����?�G��)Xf`ܖ�t�޽�J}���7�ȏT�EbӬ���M�N��yKW7��TL.�~��
s�q�}� J!�������ڠ�j�R2rr�y�jM������):ﰄ��4�1������`ꨬ��L��fY�l�RB�
�����
��qY`X.e����E=i�wXټe��m��],{zC��Ĭcc�00L���'��Ӝ�6�^&_��f��ݔ�b���܍s�4�%@��=��jq�b�`�)=S"��Q���\*^ɷ�F\]q���.��6�@�����hM�{�W@S+je~.�$��x� `�Ҫ���L���V�d�K��oiE8	�����2l~���ۿ��� �Hd���;�:�7i��Tr¿�;���]:�yE0�h<�I]H��1Z�π�S����Q��i	����FEf��$�
M$�ae��j��UGo�9�L��>UX��K��	�`��{ޙҟ�̻
o��)7{�	 ���Q��	ҹ�wO�᷈�cX /C^���jE��|��S�O�%Z��Q�a˕�FPј
ټ(��O�L4Z���e �O��?>�n sa�L�-�#UA���gZ��Q�eW�ȿ�9�5U]Ux(��,�������|�Q5-��ey7O�D������ �V|>^6j�����%bqv��Ǖnh4/☟�e�_끀0+���+�k�������TSt*���h�Ĥ;����AW_�+�&i��8ԁs�]|o}O���쉳o	�r��gN�&-!��F�!~��N�rZ�j��~h,$iՀ�{h�h'SI@���<����sMz-ٓ�'�ȇ*�IiTZqYD�l4�����}����Y�B\0j��Z%�vk�)�UMv�ůxW��w�c��v{b8���+�2�r?��et��3�����$-A���H�= ���`��.�#5�%�ه�$f��A��KXud57�\B��)��xF�����#�������J�B�!���~���3���b]����^3"%[��H#>CU�k�ŨNoRm7����"�F>�����JhlrJP�!�Ѫ;������^ ߬�kJ�R�W���#L�����o#$�V�gī�.���ݬ��ų��@����O,A%�ۃЗ��|���[n��}t�=�#.W�r۳WW��Ċ6���&3����
;�IP��J-� wK߆��u�w�hn�Y^�4 �?&W�H��e���5BB,^C	�ٺ�}33�W��������R��:��I���B�����,bg?�M^��;�O���'k�������d�DH�>l�.��1'�sQl��	U���G�rxQ���܂"E�n�+.����m����Çw7?p��$(�(���Ú|o^��Ha�,�^9��"G��ɜl���������Y��!�]ylbwu����5����/��I�Zk���ߧ��y%u};�_��e�%��b�&Ϧ2ٶ�(���s��@��aLB M'E�N�8C,{���D*�k�.2���w�$?5�b�PV���7y�=�F���;0:F�yzt�Q���~2/!+y���{�)����x��&R\��.��"[�8�AN����[�4]z�L����R�49|�Ӟ����H��FW�7U��ާ�$)�vC�Ky{����[�g�D�>�D���i� �.@!���fx^�v�%m?�����JؕQ���wt�0_wc�&�l�z��B�}�N�����P�r�؜��>�]j��@&����l�c�/o Mx&����{���ݑ~�{~w�d��*^�1�wJs�������${bt�6�fV�fu�}<2:��1�[�~�ҹ�(-�H-�K�:�9���S��9� ���z�o"|���J���\�����/L{�iX�b�[�� r�tXV�w���xiɐ�$�����C^�
��Uu�j(M")fq�o�׫}l�)�t��wS��I��;?�y�,��/J�^�d�H'W�"�~���� �{~V�a���*lն�[.�O���H�>���
����#c����i4�4:D�aj�"黡(��$��Q��1��ai��1���L�V�s`g6����t$"]]��'�Yxm�A��<7�I�Ps)��'-���vO�I�2�-�4=��6ݦ��	�����	��KƦ�X�'E�%_X��s����B�R�Q;K���B��a{�Y*��5�H	���̱�,����7�H��w�~ؕV�t�G�p;�E����ۭx �fU�v0$�e�����$Ͼ�U��"�~{�Z��	��+�\�<F5h�8�{���=~�-��ݯ��}E����ǿ� Pp�M6�'{�ևT���x�VR{4�0�\�;�C��!5ݑ�����!I A�І���\&_�,��
@F��oC$d�&�-D�N���]�cCa���n�6J���n��i�'�=�:idH�VDS�3H����+�ڥ�1�<��t1��zz���
+�;K�~�*�R��o�FcQC��l��ho����}����b�kt %ޘd�M��j��c�3 ��JFLm�5
��Gt���@"��C����W�DK{����u���p��lT��vӒ�8>qC� ���F�]֜�:�ް�]A���¹k�8T#M�Ȍ�˘�횎K�j��7��w\W�^Q?x#]�\�8{O0���F����\&�u3������]˧��n�~
̀����dL�C8��"S9����!������:Tߵ%9s�������Z:�<t�Ȫt62ߚ��J���CB�+W��ll�h|Y#.Mf�`�7\���I���z������	&�� P�B��	u�t�˜�*��ofD����/7�+�Yb�#Zr\fw%�w�;b&Ts���1FF��~.$"���!���-���|l&����dGT���+O���+H]�[���'�<�q5ţdOU�B]��(9Z�o�{G1C����+�i2��4y~�K:�'�?>7geu����2Q��E��4�_.\����@��eih5����(0�"'��(���%�2��|��mC� #�QSy�!�&N9%V��o6�o���·�{$�$ N��|nJ��1Ls����g����v�Zm0�Vy2ݣ�i����3v��] �ld�Ko{���'�� �?�U�4.Q�-�I�5���="���H^2�[|{�0�_|�xE4W/��t��L�N��z�8��SrlO|Z�׍���mљ�}���m`7�'�Ϝ��Z�o���YmK���A�����X6�aƋ)mn�Շ~�h/�!��S&Aie|l� �Y��c�y��d�Mh-�����/��§�U'��&)��c}�|(����j�Udo�m�������$�7�!��U��5D�_(Ŵb����U!��/O�HWI�3�pb�!G`�I�w�lKeϿ�'>���Dc�
�J�/ҿ�p!	�A������z���N�� �9+��e�`+Mh����V3"�pkt��P��ٴ�dx�q�u� ,2��@�p���w���+ɍ��6w�p|��tL�R�4	B� ���°��2v��I�,Y�}Q5����1	h��)0T�袂�o��9���k�Uޙ�5/��Qsq��[�J�6��2"FD�xڞ��k��_�T��84c��^�>Y��3>���e�����?�Mޕ�.v"��Ƃ�H������ �K��y]ChMXq�:ᔝ-�^�g,_�ɋ1�/3O�m"9~(o��X��Q��q�gzaT"���Z{��|x{8�VD�:*��*M�υ9^ょ�ףb�	����#��`����Iʙ3;�g���DV`)|��"7�u&�.Av��Z��]�}M��䌷.�x�įh!a޳p�"��W��(�WݞNm�� �(c�
5�����$��-\~!���w96� R�Rb�,�ǫ��'��\[-ꨚsԵ��m���e�SbÑ��)���!�9S`��t7��Ɇ���<��V'æ!���	u���x2��Ȓ. vȽ�N3ql�6O�A�Jݩ�����5L�m���;vQ?�5|⎤��3����6�6pz���M�W�x�t��u1ߗs�o�����ٹ/�D#�.,��n�,��[m�?�NLd%����v��<����X���~�s§�t;M(+W.Щ�q)y������J34�QE--�s8���u���j�~4O�T�m½�y9�b��[�7���(h��`�%�����P;-��gIt^�$Ө�a�a��!A-�V�M~��^�������V�IbT��HKQ��m�>d��ա�^����n�.�����N5������r�W�h_��<��� �~�� L
��<:a��Mn`�56r־f�<��ؼAU���$�#�MM�c-��.76�'�M���r4!�����`YUP���uI*�q��B
� �J(6��Q�>`��)I�:�<���6��El�ْT�F6	/5.gu�-�3� �)i�9�9���]�mRV��j��`�OC��Wr�����"���Pj�i�]�����kh���#Ur�����JC�ĺ+q���Ab��_�����D� �Z�S��~����'�h�痞�Oq�&?yS��!�E�<�_���w�l^|��f:�A��n�o����X@�n�������y-ꋩ$���Q�~ �o�X��ǩ��c�1kј�I"RX���%��ԍ��%�[�C.Yϓ���k�E�A��^�o�1�3G�G~��Oi0պ~f��\@�8�>b�0A���E������D����̓ATi��Ŵ�b����������K�5#�8i��j��-:v�X%Zt^E�tE2TɊ�D��?!2d�gwO�5ՑK����D���YS��Bm]�QFSF���GD2�����9�=Kk��p��/� �T��ǣ���f���"���7Ϡ���T�3�̱�/��ō�?���m�d1����k,G�,��u�AMmS��M���vdYb��>���u�1����E|%'������j����e�C)��oc�@��'y�<1-��b	�K�� Å8�4٭�P�v`�f��${l�<��H�,,_z>V���	�, �n%n�	Й��9��;�]A��Oh�i�~U��(���ja[5� p��邲�w@�ܖ���b�6��@�ha��<�]д�ŻVB)���+H�fa�L��(Z)�s��P�?m��@�92Z!u�@q����w@�UH��}1j�n?16�uD�o�������G�ɛ�����b��魼(%��
3|+;Duf��P�u�[��yˊ����d7��-\^�w�8�����
@����+%15Vs��/BΛ�$	���dy�k��C�D����Vx(�\Dh|�2s��t��c��)7�N��q�WR:��C�M��dD昆!��s3���ɯ/��������)%��*���eE�w��:1~svw���S{�O�`X[�C
��s+��Ռ���'#�X����q1�����÷�Pdb�H�$��昽�DD	��[�}^j��l~!_�"͐`^�A�b���\V^ë��'��;�\�{Lv	��}̲�=�oo5�|�U�9#����N�PAW!"����Io�c
:�9�6���0B����G�6��q
�C^����Ӌ��ģ\B�Fe��*�_�ئu � 1�G /�B���ld[�b
���� m�Z�"�Y>��D������ۯ/"�j`�Tg�+��3Ҟ���������/��Y���Mh�ɩ�1F�v�
xp`��U�Ul3��7`��CN�����o������C����^yk: �l�� !���g&�QB�7j=m��II6y�����a#��5*#
���2��Wܘ��J�%9G�
q��}���P��@�e��5J���
H��{`�М��j����$��I��V�������IFYk9e_���܏����:���"��-�>��~�K¯��^� ��kd���,rNz�xEz�}�V3�s���z?��8b@�_��	3���gR`t�SL�O�Ȱ�s���D%���zA_x�H�ڷ�l���j�KKE���|�=tp�FB9D��ih!vhr0t��>B��,�`WݎY�vF\ez��e�K�J�p���I�`*�� E�Xn�~�B�kn\0>-��>
�RZv��r��·&�`X�l���P��A+��8�k��\���^�������8��l��������N�N⾤��/�1+Qt��+f�	�{CБ%�ņce���:����c������ ]b���,�T~��Na�e�w��ܣc� ��2K�V}�#�C0$X���q��!�|�I�A�YU��	�����%u��>��tn�nf���G�q��s�,��faS��K��M�Y���4Aő-���C-�؄h�aG���ʳ f�?�URd�0^T�:�!��Ik/��x㭲�p�A�+.���kp�Z�ӻ1��G�낲M�_���x�Ý��d�
ߋz��j�":0� �&2Pd`w+�B���੉��|z������Y ?A�m{��Q���9�����e�.%�0G�.�8˘��"r���~�V�; Le�1��z�|�t�{�S*�u���(:] �q��+��	_5�<�����P���l�{��+��o�L�!E�ݳ�*�g�8�}�m��,r��8�A�ԾNj��a��{JȘ�V(�]QWi��
�Rg�;�}��p��ϭ �=��&�n�����^�r &�K�n�W�1'�lz��W/������p�r��ͦ�e̶�
2���,_����ڊ�C:\fx���2"�GALTF�(�6E!!��ُ�z���Z�?�����%������a���p�������~-kE$���>,!����9ѝD��7��5�;�b�8���U��3&6Hjq���5�t*��#��Ú Ij%J(h��g��A����^g-Bj�7LU��A�U�w�;w/5�\�RH�Xu����up1�ȿ����x���ژ�Z�-ƽU��J��f:��L�G���E�
?~�x����7\��!c^pXv::�b�g;�&U� (�vnB�f6�&C���*N�H��e1V�Uo���gîA��S<�����G�o#C�X���H��x<�;�=Zr�8���ғ��	KY+�������M8%U6T���sxRJ?\V�E}`���Y��X
2%	<޳�;���M�%�&�+�Q�}�R ��@]�H����dd�֛��&"��-+]33����j������!�nב�����vDa6Hk���3u��������R����{ʉ���N��A�d�׼m�����W���DM��]%��+�*� P���n�05Jy�ۨ9ǋHJ�"��·�ė%?]� c:^�����@X�[&;�����e�זRJ��u�h;�mݔZ�R%�~%!i[XqJ���z �cB�~0�5�P�܏h�gϘpcњ���ž��nNz$�c��C��ɭC���p���LR��\@��uy�kLa0'F{��*���*Q�6���R[S:�� fÞ��^[/QFqr�ߝ�j����6�������,���r/FP#�f��㫠�ܜN�5|�[���_�i���Ĝ�I��@5��r�ާ���|��,�M�2�V�8�@��	?��cp�9�&<�����;V��N7�n-�}��Y�/��E)��lob�X��:\�d�.�*D����~ظ)2:������5f�k�BU"a���9�̀����X�(Æ웽>�3F~��5< w��@p�|���T���-��K��P���&d��M|�h÷e�?�a�0��?p�쿳�6�w2MĴ���d���Aɝ�ډ���hC/{`� �Nu'���X���k�w���	�
�F:��u�b+���kj��2]n�j��f(ɦ��Y��������>[z���>,Ɂ��_�NOЮ;�m���E��>=V�N�Q�)��&0���KI=��Q��z��{P0NaS�n���8��?%�QK��_���&����m�埐�-���>�C4�ki�@-H.}p�-��#NO3$c(Ba�����,lz�4������j�Ɖ��kElwV����b#T�rM��k�pF9:��`Y��G���XuJ��0�!7d�e�gߊGj� ˈ�H|�
�\�hf����o����XM1y�X����+զ&��"����z���ά�d����ZQj��ڲ;gc*E8�q�Ѻ+0� �kQ�B�'? UqH�C��������p1Я����eK��k?J�"碌�ѓ�g!�r̢W��g#B^�3=��2�v�b,�Ҩ�2�_6a̚y�
3@�m3�9x[5�!�@��.� oL��S��{�-H�6-��~K7���A�8 �wq�,�����F%�ĩF��X*����ʘ��z�y@'=Vq���x���&H[#`n��ch9%�]dj=~��ag��J��S7�Jc�c���j������mI�-n�B�j�U, �Z5^������7�Zu�Ň}[���y�5!���#����׎r8Q�z!ǻ	�^،��:p$T�aO"�Ԏ2�C}<���\��X�0 Q�bP�2Nf�ۥ�4��S�c��16�{�-7@�Ca�>�Y2(�T�t�<��,��b��nHc]��=���ɪ�����Y��8�u����t��q�]X3�k�(�߯e���
�{����7Y�|��5K�0�<�Y������Q������g�`��%����Z������<Y������p�7E'l���'Ƹ�OHpvd<:�I����q�p�i�W~5ހ����9yr��H�)�)q> �U�^2��zK��o�@�3����N��X7);�
rC�(����Ù��E.��K�i3����7�oy"Q�CR�si�/���k�M"3h .P�gD;�����q�Hh�^�snH}��1&f�I�τ���K�����9��=��C((j��NF$���{ �����AM���e�p����ݡ�*bC�@л@$�Gci�m���
J��#-�H���I9��H� �|dF"��m%^8?xA����7�bx��*T=�y�3 �A[��pڲ��@����1D㦾�3O���.�6�`	#�NU�ʳ�˖��d�H�T�<R��>��%�)f�M��ð�8�G�9�q:&3;bZ��*!��Ż��葟�y�;~���4����O���]���37/o?�?�øݼ�f[���]tW(�d�d���Ͱ��jSW9�����X�L#GU���LhŨ��b�.�LͻM�Ҍ�V{@y:�*f��{���z�����-@6��ano�v1 ϴ�:Åo��< ��kK�Vve%���h%��kC�ndU��a͌88��D�cyOQ�H��$L�)v(��]��-���cNt�/�дh�0A�<-����Ǖ2�Hd�Y�C�\��[�CZ�����!�ld���6s�Vڸ��z��jdx���F�y��Lؓ r�]A�5��hd��Aɼ��7�E1�r3Np�!��z������?-)�Ah&Űdr��6�)��5��� �h*��c|G��8F���6�}��Ă`ݦ�7������X64'��"M���:T��F$4.�,�B���ja%��[uB+����pU�[��\�-��/f�����:Zْ��u���ѭ�jdz��5�t,��u~�ZM3��E�\��.|�3Zcj�K9��VM���G���O��t�YV���T��Zf��9rg]����;��/ �ys�Z�!1�R�;�״�����A���
�%W_fx�A�r�zG���W�9u���3�?;[:��EE�>/�恤�(G�&T ���b����lg�)�r<.��p� 8*g�Y�ςK��8MNўB8K���w;�;}ϋ���6__~@Mj�>���CJy�X�<�̤(~��)��Pal�.��XJ~|�'��Iʿ{��M��Yd�︱p�D-���'��8T�:d�KDuD- $q֣Q]�U��W-շ�@TC\�g���<"�J5/��C�D�oK/���H�b�94E���7��ZpKc�mf���#�ђ�6	�D��	F��(�Kp��˼���y'�7듟��f�4s^�����R
����_>�h,+�qo�3xn�|;��V���4���L������rV>Ѭ��_/ �X1;`�35�$���s��7�*{���I��i�z�cpJ�~9AAO�����)���7u
Kx��&�Գ��J��[��K��(Zsz��w�.Na�l�:J�E�dV�P"!���F��}uͅk���$t*<돀˔�6�RݽU�C\e�����V�G�N� %�/�ؽ�B|N*:�q���>�{��A�ݦB/DhY%�z���z�wp/�-QE"����鐲����?�6BR�vg�Gw���~ydp������>�N�X*���iS},��IG���xkl6c�ʩn�ʶED�8*�bc�ȑ����̎�K�i�O�X���j�T<2��.lQW���!��	-qj���i��Se�1�����v�4T����k2�8Zi,Ew�N�-�B�X��ѾOh�VVBS�^{Ƒ�@�o�X�}��C�3 ��ȵ��6���ia �ԟ<���;�ՄV3oa�y�@�Fa��^�8B�@�T�6�'����Ќ�UA��=W�"�Bߧ���iyd.�\�
[;'��(1Èh�
�{o�
���Z���z��Xu��6iV�Ǣ򊪳k���[������s.!"��A����`o��8w�ԺI�صA��C�h�Z~��Ȩg�#h��*BE���4��K�v��'
n��}�%���y��_��l�2�n�,�
	X�%P�9�=�Y�L�u�U꾹Fh�S|͈톧Tm�q������>X�E�a�m%��99/惛�Ʈ���+̫�{�=�福��U��͏��wad�	�W��^�R�/�R+VY�n�c��Ľ���0D�����MO6׽�1lyZy,$=,q��.��p�������z,o��>{V}9p�K�%�9��퐂^#v�E\X���9s߹&��5����
�Q��̓�~�M���#�Ym#K�g�d�f�GR�r� �(���<��+ k�X�V�Q�I�+�1:rm���֜�7�ݥRx��X�,�������G�������� ʥ����[��K�$��l�:ìhL(�-Z�ȇ�UT��I��@�Yd'&��R:�{����)홋1*ʛ���T.	��U�>�N����:����	��#��n��U�Q*z`���\�-¯���k��w"X\1���/�uK�Ӏ�_\d�������Gk�U0�m��qL�0dM�L\0��T�����p�~���e��fS��f`����_����Q�b�`���g[T�A�9�t��IM鼉=�(o�mP�O�@t3E&}���E+i8D.�F�g���Tf{��Z�ς�?L��Q����ף�@�k��I��p����1{�g�� ��#��?g]9({��ƭ�'Gߠ�_?�좎�g�ue�V�֞J]�Q�3�_Gh��(/�� ��0.<���+;牸�(qxs�&����KQ"H�{<ywݽ�X��$� ���Q�V���"����a�_1�{41b^F_N��G\��x��3-,I���"C'_�˘q��؟XjD�`���F�v�$U3ou�d�(e��h&��\�,e!����%[�z���YQF6H�g5"M��Ǎ-��wQ�i����{D؄�X���Db�����N���T�q�.M��:Ї5?��n�vy$�8�r��t��!�
$���"�7�\\U��q��'���d���J�!N�.���ח��ZРA@��P=������ݕ
�3h�F�z&�7nQ��	 �����+L�^��`R�{���`&�UG�
�.v�/�sѥ)TRP�.\�xY{�+>7���͒闉�<{����ˋ��/,D��D3���sa�K�kp��%��#h,]�4i��jq�Y ��7��t �h�x1�u�o���K0�J��-��v�M��= Z^*H�֏�4�6���9X^����� �cH?�U��K�Ve�Y �n��`�W41��5O0�?�^��V��o�\�g�IO\�'�g���7ݙ��lO�t�ص����n$9�l��U�>���y;'�+�a�h�
���;6�vS�0�:!��fট������-�'��|���ٻ-
9;֏���T�#�򨤳�ؔO�8��%�)g����S��DʹT�?�[`� �<�C$�^���>���n�?H�}���(��q �I����9���y'�{��]�V����ӥz�J�uG�5N�߄�w������xs�{�����I;���M�\&�(��=?3�Mњ$��y㻟�ѫy0Y�ݻ�cV'��9S͙)����aYra�O�tA@�z���<��tT�'K���C	���,�Thh��nVx��Ԕ�!��=Ue�-:��e7�r�lJ _�e�os]��`�r��������d�E����N
���|܁����4:ALPYoo��;	�����3k�>��R���E� �s<� �mMOh���r(ʷk(��?,�+!?$��8��(=��%�p�^Y8��Ll��Q��e�sy������x:�O�fQ��ֵ��ă�<a�+-���T�T�~w�ʌd���UA�Oh.��P8��=������߱�d.��d��(����{�]<d���R\��"XJkU�,�e�܄}�/�7����Og|O�4���A��5቏$.�#�'2}�duY ���'�[}�}C(�(F#/a~��%�5���k�l'j�����@%Ғ��8�.3i'������I�7*�)��ɐ�;A:s
6���������@�]���"_�<q���=']xo�"�!e�-h#����i;�y5�Ѻj��>�j��P�:���ʛ*N:UD��&lk�Z1U�����ф$���%"��Y�箧O��<��
��$Ш� �mR#:�iف.,!��t���^��.�;�d�fN�?� lu��zz��������a�H]� Lt���N{Ğ�=��1O����8M �C7>�h>����-v�,s9[
�;�t�D����^���Kf:��z�-j��L"䴺�ir8���m���6��B�Jiȥ�Ȋ{p�}�U$�_�/����j)b����2��yb�A4c={��
�ͯ_����xL	(��� l��*i�����f?0��w�/��6�&����Ьƙ�p@!�Œ&��}����l�JE]mh/n[i�ծ�C���r�]]�qJg,_%���h�GxV�0�����/�&(2{��� ���[��(�L%�fK;�LS�T�z��>/�L:�����P������MÕT�˄%q�W`q�h���M��|����=��!��b����q��.H��j?�I`#�:n�%ю�>�h���Bdܡ?NŃo��e }�H6��Õl�T�#ShȡAH���<�U9s�=Z��L?!��iP�$�pXB�bHN�Xvxku@���C-�r������* L�5tC>\���͙�C��ﷴ��tv���V�^��2�9�TȽԸƔuu� �����4g#���U����5�y��7�������J6�9����v�?�l·�>��qǥ;��E���c���H�����x0��]v5yctu<1�lc��+�ʺ���`�2,y�ϥ̂�>q5��4c�:�+i���dú�v�;��q[Q�����ɾ����0}	�P�u�y�;�01�VX�n�����΃x�)8�e�v(�4�ODJ���Tb����'�5��N��"���,� �H������O�;ҿ�N���Xy�S�'�����j�o��/��=s�$?��
��\�V*[�7_^5ӈ���`睎L9�4K��Xv�V�sg
f��L��4����^	�$����]j��lb�J?�����Yud�s�$�|�J�Ͳ��s��S
7T�����w�f��Y�3eP(���3w3�&K:q	C.�c��C�Iu�Wجv�Ǚ����@[��"u��a�WcX�m���0�>��Mm���N"a�{����mu���O`eA���P�y��<p�cE�;�����Z�NI*u]h�s�1� {u	�U�޶��R���u�=QLJԪE?��kTMCX)�/��ۍ��c���sJ�oq0ċ��	o��g`�ËT��~���ם�����ձ˼7�߿&D��1�9	�K�W��έ��F�����d�T�;z:d���<�V��H�sJ�Þ�2q��BT�5rff!�M5����݂���,$����+x�j�e���e������Cb�S��1Ķ�5��?Fp-�`��4nF��������P�G!�:4��۠�:��$!k�=]��}�c����X.���g{E���8;�ؿ�[͊�F�NW����I^��]�&������޸�F��f��A(��ܲM��?�q������6{��8��k��좽�Y���e^�A��R=2� ��l�Y`���>���@'g{L1IT�@1\�烃��� ��O(˚�1#k!��t*/�A�w�(������e��9po�O�`E����ٽ6�&Ԟ>�*y'��L(�o����Ұ�j���#��C�1Ow���JQ��\�OZ�oq�q�$O��;�Wv�� S�+X��N�U~���:.*L�o�G�\lIy�sy�4@�T�$�>��%��E�:Zi �
�c����B�U�`ob�^葩 �w��t~��K�4�Ej�qj�~��{�B<G�!�b�( aTݞ��x��>f�;��������'�e;��ٖ��n���<��)y$I�H�4��o���4|��D�����!��E����m�P<%(s�TsřȼcDe㰀 �m~��9���4o�� ͆�b��:y&�T�/����cxbV��7ˍ1�M�E$�n���f���x��9�(5��Z��i�rN�Z�87So���	&V*T�ߤQT�	�[�Sk࿉K���C ��1o	���oy�P�߱�Z1ڵ?��}�A{�R�ho]��*�g���S-|Cv�f:�''ʴ��(�k_���T��ӆ&.�b��n��A��C��X�41�+Y8�!�(���0Y{|h0' ye#��=�gQ=z��S���vΫ���)����k-39m`y��p��4��eo*R6���O�Е���7�霘�t5�'*>���P������_es�.�݅����{��[��[��y>� ��(��2m�>���HKx��;�b��o�o�6�1_	�f�^1! 8�|N�zY��i8 /�`LDi�����N E+|z5�4��~�!A)�Z��6���ߞ$m�4%�95�y~�0�W�ZGF!�b���1[[�g�rBf��M�ZQ4P�����=���� 6g��W����%	Bf��;�C�d�G9x(��3�'������>"�=I���\Ԩi�-��3��1�M���\��r�7�(�;��cj������ |��s���a��,�W�jiD��<�7R�u���+��q��B3�"�j1#}_�XLd$��O�<�a�jh�#���_�Ujd,�녹k �x]�bE|��x�	Pp#�a��C�*q�̞������Cund�ݒr{��ؑ�@6i���	���*���D�_�lS���s�n�Z��E���0�Q�'�Vδ�Y���ozo����D} j�W�τ��l6�,Tnjwތ�{��-��mL��Y��Ǧ��iRSn9���!��R��)N}�~Q�C場�{C/�,��
hYt���;�����yd�4����]����0°��[�<�sq��\B�g�B1�v(�7ߊ��\!O0�]���� -�n�)W�����[�������gO�*��ښ�g��Us7�oi�d��tS�Jx`����9��[���^f�O�>�c������G�R�2\ćEp�>�2D�����,4�Q�� ��<��zNG����af�N���E,k�Et�H_���檊VT >dhhnvdRC�:���mFO�������|�<o�Ĵ� e�՞K�GT�"!i�Y!%��]|���AYJ�){B�2�Mr�[�V;���{������<2��Տ"��{�K��p�<g��pݪ��t�Ͳ  ���rl�Y u�aY�w���8�v6�����&�W)B"m˾-%9�^��3}G�tH��;[��w����� ��1�X�������|Тǲ��1��V���z�!g�ƪ4&'Bֱ�|�F���
)����%����0&���]�6��+b��*L�[�A����u��y��̻���V��6��u!׉}U�K�S^3��ؤ�+���]�/x�3m}-�)��������H7,�j��08�jV� ��-6x��J <~�V {�A' �6�ɻQX����`G�>�_�up �2����	����;QΕ*n����$���T)|�k�NoD9��V���:�u|��9��Y�H}W���t3��T�=];��T�����.1Ym��?(�(�f(%������O'���땝|���ƈ,:Ʉ�\�5��9O`�ͧ��ɉ�qaO�wxG>�fxt�0b�^wlԺR|�?br�&�,9�����(�?'Y�n#;ca(8��eR���Z)"�G��7�W �C�4I��OR��g� "�$��=��kuj��b��/�����::;�Bq��J��&T�x��}�� $ZЊ�L�d��{�4��]���
���pD ��]�1�?>TAY�;���0��x�"�6�
[�@/��UHw�w��?AD|���*�t��������KV����.!�ȭķ���_��!�9����?p��
x:���W`�%�����$A^�\L��q�=�w�+�v�'w�)}!)s����t�#����x�X��!�^ T��	�79�.����\t`R���D�,�?f�%J�����G��]X2����`�m�)���;ۿ�ָF����l�������$;߰�jg�6PFɳ��W��}Pz�N7ySD���_x���Mf�Uiv�],�vعQ*��'cI'X�_�n{ч�4���+����bd��"E�w��]T=�tr&,���Z]���Y;�=6�V��n��=o,����'��.����i��`2��^z�b�_���S��W���3Ad;��X��y�+.ŰJT&��bA'_#J"����oi�8D������u�$�$�$��M,"==�{������J^��u�O��
�z_�a봸w�MKP����s��� {j:,|���"	���K;{\�o�L�*I���=W�Ө���#��j�e��圀>I�5�<�����}]��FM��Y-�E�X86�a���(�Ґ2-��і�	����'	A%{;A��ǫ7���2�b%u�]�.���%Ww����u�NR�v�@�m����f�8��'cS`>y{�:ը��f�"�����¦�<��UA����IzT*E��=F��:E��vr~$>@��v].v6����J_��:3�2�M�̆-u$Z��6ݓ��$�T����4�C����J5@���!���v��:�����f#�6W�	��*��N!��K����W��7�GTY-AY��F��}�i��5B���mT��DlI�ʅE�J��}�Y<�b�(bD�x�����pa�klճ�n�A�b�#����W�0��1����<qx��^S1A��^mI�i�y�"���B��3N�&U+��/Ev�ݠ�o��%�r�u#�s��1?��K���*;,!�� �H��h�4p^�:W�M�̪İ��dʹ�d	��r�)�H��	��-��[�G����%͹@���()xϏ7��r�Ѹ�2���b�Y��� ����~��g;tۡ�S��T����W����6J�� ��6�.9�?�	����Q��c�R�I�컞V�R�]Co%�$����� H��*��H�����x�ڕ/]:N\�y�sI�w)���y�w�3	4��/claŖӶF�uP�'
��ƕ8ͻ�팥~�0�*(�C���'�­w<��������$��+(�����8k���ݷup���ҟ`�Ԍ�� Yø+<��`���TwͲ�7\�n��r�e��}vV�G���_V�;�J6l�����4і��q�{�G�ua_`�<|Gj�مk�:~~��D����Px�Y7yE���M�UT�qL�4:A��jq�[�|W�o{�@h�=��� � ��Z&k���j1���_y�ޒ���D'�ВPm�>;��yd[��ە����7�V��h��5e�{��4t�cv[�����n�J�Q
Mq4�:	|*N�jQ�H�K��� �r:�H) �Z��ᥟ,k�'q�����^�Ĺ����\��L��)�)��r��g8ƠP��)�mrj��`5B&f\�e�k��P-��b�圕t�<��N,������S�YM�9�l\��X�yQ�[Wh�mmL5b����l���Pf{P#���f!��f���PKu͎|_1��YM�17�[z��&��.�,Sq�T)a��WD��vH�^���4����
��@~�kǙ�y��A�^��SĞξ�򅟨w�*Q�T@��E1O�p@p�.�^�㫠�l����PĚ_㕍����\>*"	��W���W�t�k(�s�!�ķ����'�n���ӫ�ńG�v����5�vC�����~�]Ǩ9����2��9�B�"	şD*c��M>���v��ڿV���Ӫ<o臓"ʍ"�s��P/:��v�J
�3��.y�V,xxb�/�]��sΧGm"٭G�{�"�J 0h���y��n�I
G��C�"�F��e�S��D��� t_��/�N�����f�� �+/�m2����3	Pj�^�o��Aȑ�td�\ �A�����=[
m��+�1�YB���W�i|�hV��������ߞ"+lt�!�ʨsG��+�深G�GF��K�I��V;������7dS�����}e�ߓ叒�j�;O�l�C�_�����U_$��w(�堕� kc5/�]��тN�h��j�DJ_$7%J�K�8Ob�D�����x'j�T�O�Y��C`�� Z '<�'J��\���'._瑪oJ(aJή���k4�5��f
�2� 8�#�x��:��z��Yn}��7��x�?5m�Y��L�&�?�W �:Y9����4t��!k�q|p:��"�Of�y�Pg��a2x��0�A�+yl��Ǉ�t)���D@_�8H�=$<OeWO��y�;�H�a��S�V���L���n�����W�<��6W�XE�8�WG��O�}^.��q��/���Ö�6h-&'�4�V����p��b���5��>���\��[<ӝEd;��ӝ� ,ơI'�X�H?~�sK�iN(�+���Z�L�[yu��c�u7�.�چk��+����xԶ�/Ϝ�J1�'4҂�{�"���#I'��I(�".����ԓ��72 A�������x���ӻ��C,ٌ�0:/I�,�Ӫ�@�sK�Oژ� d�A���Tk-�U��82D~v�
�/��[��.N�sj�A򌶁�q�D�Z���@(�It�Y8��i=�X�#2��?E�٨���['7/e��"S���)�xYw�I�7�O5V;P;w���N���?� ��7PP�����Xk���z�����˔�٥d��_kG��7���2>0m�$�b��}D�G=�����E�%]�?p���{�q�ŀ�w����O\TJ�4⼱ek�sƹ�Cw���C��pE].�3/���^�!�O�W��t/Pph��ǣ����q�+�E����Q�<nJ2�돻�ĸn{�J���e�f�c����3�����U��#�yb����N��lQ���f}g��S�١&�1*J��;ts��N��ɩ�>}T^��X�4pҍ?�E\ݏbr�z�G��cV+_/;�ў�Q����=�ǹ��F��羋�Y��c\�L]�$qc0����ݨ�,�7��n��#�!�� ���Jh3�wGa������1V�=V� �L|j��%�(Gs���vM�;g�-����o!��g+�&~�Ov-�0�ˈ��?1��R@�я=�**!���W�u�߹���	 �EҾ$�Z;�n��O������LW��7[�Yb+��J��
`�?�z���b�}��/��rE~{�9F�G׾ʄ�ބ��&�@>��:Lݪe���o�7,.�;�=~��"�t����t+
�5D��E�+�k��[�c�h{䇓")�?3w��*���K\�0Ka��g*�:������a>� �I���ON�?Ù����#���W�ֽB`�����ܕ�=8�SӐ��V҂�g����#1o�������(�*�=�����d9{w�`��������ǆ�80w�=c\ ��F��D��zL���
�|�R,�'/�N�X��o�D�U^�s�+(�Y ���\Du@VQ�!�[(��&��dݭ-e�>���	���3%�h�����I":n�l���N:�Uj헦8ڕ�F��K��^6v�f�0�� ��ԩ���L�&�w���Ȳ��🙘f���u��RV�
��:Z)�H� ����(ɣ�u��v/��%���d	:�~-AAkO��	�.�6�/yW2ȧ���ߓ5�d�jj�/s�2��/�ԛm>���2-bn�4Wj/��=��(F
�N:؅��Y0��|f�G�4�:D��B��r��5rNh���ҥ�u8�L��x��q�������ӫ�����<�����8�����a���YZ��u��	uFy�,�xeٶ���w�:�6� F���0Nu����LYk[�m��y=k�3j��NM�{�t]�wz��es�[;'�5U�ؕ��,uv��9�8&P_">bF'�����J�6�y�]ot�O눅sd���K��:�#u��)6��dHU{�@�K����7����ۨT^�gQ�F[!�I��b���S�/f�_��ؤ_�Mw<�SW+�ﮋ�`�x�g�#��)�iP�d��T%�n��y�1���P*8����y�ޮ�G����x�%��� �v^��z���o��o�*+&�t�oT����^�Z\N��:&�:�:f��,n�,�l�@[���`�7�|ۼA���b
���)���b��m������F��C\���>v�E0#r���렀���c�ωt��C��(O�%�V�k*�h=���͹-��z�8k�~Y$���7&�P���.�u-���N	���W�`�?(T�Z2�ݬ�<�����z��b�f�NռB]e�a�y\�4��5�5O���4�����V�������-�?X6�����b���m��y�ZG@c�Qֽ���0��~|a���+��K/sN�C����!
_� 1@�Vf1b8�A}3Gp�M�椊Y��´��w�n�����O��z�D ���"�3D��Y�F�6ڲ�|�w�bX[w����*��{�zx�ua t�X�(�wd�F�~�M��rp��vO@
%�k,h�6�5+cd��"E�h����p��I��+cҀ�%�m+ ��|5j�K���v�Ptl�%Ԩ�J��J�ǛLBu��^X1[�F�e�m�]ͻ�Zh�� $4���dxm�������I��A�n7�[�ӘI�[@=�[>z�h$���y���� "�؁�-"�Ce/�!|ۋ�c#+?Q��In��8��H&G����h�P�&��{�р�4:�PxQ��n@�F�
k�7y�z�%*y�I���}�?��]haŵS�|n\^�\��-xQ�f;�.�8D��Ïg��] ��yAib<L_@�-�|P%�I7'�ҏ����1�- �	yN�ݷhLM�ov���d�)���E���R��!p�;�6M�r�Ȓ�HW�\�����:�2E��.�)���}���:-�f{�E�=��Z�C紱�����ݕ&�n�~����'&MQ��b��k�����(G�Fe�H
sY�#����G���<e|%�fv��20}�:m���p[�)����e�&����-��a��6�0���7з$���&��4�㻉&�#~u�gV��2#�LS��:ŁV9#�,�z�^�%3b���H�6�L���λ�J�"�0��ӆ�x勓�
���
�cܙ7�E�mD�Kka%��2箎$hz��TVM��ܿ�}���*�o; Z��f�{TJK��_D&�~�o�Ph�x��uazr\�C�X�� �.jKz�U�[�dF���$��.!	�� �7�<��b��;�DN1ѥ�e�sq�'nTW5����LT׊�;	^+hI~����`lCO��=�g}��0/7ql�̬��
Z)`��|͡�mr�)QaQ���R_mv%L<A������r�W�c3����uK4eu��B��l�f���Jspٻ��nA�+��Y�1�(���Hw��X<V�Gݲ)�OG���l��������(F���W�[�0%RD5&Z�_E�~�y��
N@je�C�O e��Z�6T��,���A�����`϶��d��]3G4/P"��|��	R��⸏(��þй�a!X�:�9튌�]��<�Z�У?�x���Tʏ�n�g�-R��\ll!S���=��'����Q�����ͼ�d���@W@�	�l��(o��LM��z���?R<�E���z��o�	a^3	t�ai$~4��!2Dċ��U��d*�ʬ}m���-V���lMK�Kx~�N���w�ۜxV|[�n���Pa��$��*��>B�,�a��o��ϔ4ݟvD��T^8��H+wb��.�k��bE#���%��B ��?�ЛH��hj�Y_�T�Lnѯ���|@����?��;��ṭ �a	���z���{%�D��I�b���O�%���CQi���c?�T�_�9H�ߙ��f��B���yl&������W�l�����0����GH��|��1�C��?'����o���^?�+���"kGo7��T�x�Y��y�?��WnV���B>�����)R�/!ҧߎ~�{����o�ݨ62��D��r^��M##�P�BBU��AOh��"�pl�y}�ǻ���Ѭ`Ω
�������;��K��l��z�U�.�������,ɼ�|Q7wG�_�1�_o؈W˹d4`����7��Rj��S ���+ӋVT	�0�YM�OI��ϝa��	S�n��K�L�T�W�5|�f%����گ���>��z\��{�|,�;�t�)��� ������!���|��h&��������'�+�p��f�ґ�:L�xw�k�͐���"�	0a��]s/�2ʲ(���e	�����	R"?�Eu ir����n���S�N�̱�IR&��^\�U~-�2Rr a>�k^��É)���>2����ɦ�6g@���Ce&��I���z�w�x�'�<�
�R�����	�N��K������yjFR瓬9#.�D?�/Kj 0��7����^HQhO���&$$,i�����1E��&(����j�S_�ߟ	�I&#��6�=�8�#9��?A�n���:T^�!dt}F��D��|���PW�`W	��[��KR��c�vr7�|}Ǌ�\&�U^��Ƕ���S�T�&M��그�����I���w������xk@?O�ra �(f�wB���~�������9��)1ML5X���;(89�>zI�O&��H�j��Ǟ|���!m��Zo$��ڇ�7|�g)+���]L�i'C�7�A�:����G�x�dʚ��b��ۮ�Wп�9�Bʽ����*���_��l�D��n�L*r=]�?��eHP~��+c�������%ڻ`��.#nߊ�� *���
�oҎ� �SB+��._|"2���MG�@�.�\:�����ŀ� 0�Up�#A2�=�R�N���y����~+i.GR-s��Qб1��z���Q���v��q�;#����K�/�"&��� �bB�9��8���9'S>-���n��t�੉)���0����R��N؜�9"�x�W�R��5����B*`&cLO�45�I���}}j�)a��õZ�&gE�����֔T�=�������A$JձN�H �F* �D:ӴGi[3 ���QIr�}�Gagԥ*�9�[�&�-���z�,���y�?sx�pHԿ�D����J��rf�b�_6X[�W��]�^��Pg�-z-L��)�����2�C�N�Z��+C��p#zEUm�'�kp|�L�ʙ1�|p���n����v�6��6r��s%EW��υ�\��)��~:�:��Hk�pTwExbC�u���$w��D$����%5��� ���x�ş%	Wȭ�СhME�Z���3��������-M|r !���1Kv��Ӄ�j;��QG4%�ۧӡ�%�s��5�������;���\��rK{\F0/���`��VFL�L�H��hsS�qp���uI���?ב�BB[�A��L�m�Lf�a�y�ƨX7�v ���a�>�lQ���t69��<�7���zۄh"��s���k�I׿�1�j>8�M��I�2=�+�#T�J�A���@�1a< k��а�n&F&��ߧZ��|hF�l�` �:����4���k!:�[x2�z�ʋ�������tonG�Q9�s_���.���|�|)DU�e��ma���9`���f�M�#I��O��S!:6	����jb���k�Q@b^uu�sK��|2¶��M�}eN
�p?4��,�yR�-�:��Dj��{�0@j�g!!&+�˔��2nx�ڂ/���Q7kU]�@���h��s�������Z�u���p� �r�amW��k��u�p�D�Ϋ��!W���PP���
�a5�`�����"̜�o�Nl�C-�*L.�}Ç>���c�ǀO��;�}���D������p�Y��P�؝~����	�|�Ss�P��ﲿ���t�X�yT3j�6L��7��8�a�]5��e�P5�P�CK��	�UGi��f�d�Y�.{��UWb�����b�W3%�To����0��C�!u��7�OMi\�ޞSȃ C �����_V�W �f����H�����U�%��Ei59'���71lGD�F�K��ӯ�M�o$�P_a|u�]�f�H � �K��@��N�A�e�}���e2d��F����mp�D�������E�z����W%��2SD2�\O4�G�f�� �f#.��_��1�6��b5�}z�c-k F�?��q��38�k��K�`����\��o�T�o�=V^Hi����O�Re�T�����
���f6�BƍF=��s�����{�y�:m�9WP.�iN���fҗ�s�0��b�z(D���Kޘן��ψ����e���U[���wj+�~�S2�	�괚u��)#�g�k��C?��z[��1����V��2oZ��3a4�[`�\�4[up/O������`��A9��^�>����?��3� �]j;��mt��g������Ǌoc������hv�/տ!�<BA���*T�V�|��.|�빃�\PX����{��B�����H�W:r[;Q���~<SNK+�(���߂l,�g���3�ޞ*g�)Ѥާ��%ѐ%B>�*Y��1#��a��Na�4��ha
+K�ϰ�:��ǎ{�S�D�s����qlLX�=k��B�,��PN)
r3�=֏2J�󒵻�����\ΎΓ��$����"'y#���(t�8>hd�Kqn�����#f>|~!e]�3�G�����-W�M����L���	Mi����薖����lJ�_�#�{��Y��ᙱe��Ř�n��C3����B��.^(��_�xg����n�����@<6���և��:bn�]�U�r}�[;it�?=��Yx�%R~9sn���F�X�l�0}3BU����ޡ��W� ���=�O�>9P�f��('Up��ĮPoJ�L��	��DLC�x̀}#�����:�z͡������ځ��u,c#�L�A���
]�"U�� 7����ޮ��&�U�h�ޘ��Xu3L^���yg'Mh��l�'�SK/�vJDOA��^�{v�g�*�G�:ŽnP3������������3,���"���)�T$��PM�E]���p���y3Xž9l��^��Ͼ�-4W&����)�/MB��&��\�â��w �4�J�m�\K�����I]:]R�4u�H:5�Q�țq�� -�&d�����֠��h
��f��M51w}dO;t3,\��2B��P<��O��� M�Wh�OJ��No��2�i|�E!Ý��e-A�����+��M�虚K�,M%f�q�n���^5Z��*�cu/�	�$]�rT-r��?�����8�i�B$zߊP����B���_�Đ'���|�~�ϳ���s����~�/�񅭚�Lꐇ�P������wڔ�Z�±m��8⧑Ԟ,UZ�>ݢm����.�l�#�U�]f��XN�Z�][�D�@����V5(�-��u'bCo�a����6\�8���0	��=��5���WfS�t�c�
��Ń��n jf��W]K��\�^�1�%6�l�m���͈5���-;�'�PO����M��`�d��ƣ�k��Q}�956s���t��ԃ7���ob #���s��/U��E~9h��x��s�;��`<��Q�I�k���I����%0̋�<$d��̂;����1��Թ%uы0�Jʽw9ݙx�-��+�V	�7��+�@!pF=&�#[��@�P�o\Ո�ި�����կ�A��t��{@���A�H�oH�Y^�L��|����ț�?&\�K��h�K߮�Lz)�i�ˣ+�[����J�W�x�>A�kc��w��:�I}?w�Ҧ8r�"�~aF�I#��'����1��ln�<���A|fN�j���۝+����ibX��쵟;����,�o�r�n�/�����I�DF�(�q$�Z��1��t��;hro���7�^��B)&I�|>]a���"�:2��J�?{��1L\:��&�zT��>�o��U�4=��� o����
��c�Y��_�cpg��xJ��2Y��G&���{��ށsk��i��y������Xk�ۙ�\?�O+����՜������5�4�O�xw�ڢi>�w%ڹ�p��jޥ�����u����Y��Rˠ  �����V;���ׯ��OўFF�&݋�>���zg=M}��6&2A��I����Q��a����WC���8�(�����cfL�����:�#wj��C���jЈR�D�?��q�j��I��z!��0Z9��܉}�Y�\�8팥�l���T[v�,I;f�ڨUjV+��W�h�rQ؊}6���<O�h@6`��l��#�l�������@�<�|k�Oyښ�������Q����>�9�Vwh�L�]�D�5�U�P,��w4�Ϣ��e�%�@�ޤf��$l��[���{��+p�@/Ud��@���������w��u�E���^��X?��^h�1uG0i��{*��U8*8K(4����E�)��H8<*{��3�j�d��#f}ԑ����62��R�C�ڪZi2��4�`Y+�W�>�?�
;�����l&C��2̱�m�w�>�U�wq�M���zE�X怈��qhf�H�d��O�T��f1��=x�����U��խ�Ыu�J�Y�pL[m�'�NN.�[��;"=Qч�H�Aܜ���.�?:s�KK:6V�6Y�����2ۋw�MúE����)���g<l&���deĦn�����;�hQ���<	�2x�ғT`�	�gU��9B"�=�`�@ԣ]
��?O�D��J��'�<鴂l�6���wzOB����ǩ�%��~l�_[F�xo�KF�����r�_�k;�֢�a{l���S,���1=Q>zGXnY�V�$�Wʗ4
p%�B��3�#���W��Xa��I�v�v!�]~�:O;4j��KI��"�1�d��c��.�j��-i	1���j�Q�W��A��0���솉�`�}₩���R��W�)��\	5��<��t���5�g��_b�nj�����×Qf	憴´��������Q�r�wP�[�Ⱥ�}�L��)�&;����LL$絣����og�1� u�硻C���q��?�Q#��͖C��	3���z]*�aÃ$sm�E�^����f���Eޕv\�ĉ�����|?%N
r�4�������/k<~4�����;�Գvl�+޵�XZ����������j�O�s���P5\�	�@[$^�CҐi�r�!aDa0\8��O׆�Ӗ�e���/�I��v�ě��
�Q$�CA�Q�ޟ�zEY�Kct�b�CYN���j��0��;��f��H�nh�U����0["@t���.?hq$\�M����b@��T���U��l�]�6V���Su����������} P"�a�~�Z-M�`IĆ��5�%{ �=�[���)�֙���Lb_,��i n�:��0� @PP�6�	^Ui�yw�g���1V�]���7��&:S/p@�����#
�����4�.�"f� �+�w��~��b[����i�^RCy0�%���,(3"�	=\)}�D�͸{��NHs�s|!��&�G������	B�3��b���L`���m+d�zx�a�ΕSǟ!�ʛ֛A
]���G�k��Di�A+�Pi!�)n	�S��
�����\U@���X�:&4Í���ZkӴ�J��8���
�����%$W�,%�h�{�z�;џD���ժ��C���	ލ�s�'m�Pޣ���;�,������v7V3�"�{�o��MG�A��q%��궔`��!���2(�a�L<U���$�f��ȃQ�P��ʕ�o��^�Lu-�R�����J��x�v%����J:4��M�m���U4]6��S'>|Ѫ�[�A2�*��~,�1i��-Wg�c�M��?]]��0��
�G�mf�I�7} [�y_��V�,"�.���sK���.���R�8�x1��G���
����1��oQ�Is�R}� ;h7�;Ww�m-����_�԰#�j��R����pq�Fɺ�!.��C�/?g��Ð�T|����u)sz~z��'F�z��($�`�k =�p�	�_7�1��:��VҊ߆��IT�E:��y����c�?.a��s1��ЕBu(e |���NV �� R1K)�+�1�Wn� $8��Y�dY�xGRO��߃R^�!nγ�iw�eSיf��~Y�7��#h��ؕ���6]��:���;���P�$�ig�Y�?��ЮR��=F!�ih�g0�a���M1"���ľt�^mn�cv�s�L���<H{X�߆ɨP�Z3��q�+3
�)Q�L��ݞ+�޴i})��"�@�Ā�t�٥�= "7��з�'Z�$h2ב��c���a���x�wӌ������g�T	����V�2s�=��@�GV=���6aH���V�jt�!���P���R�v��S�a��n�tt��Ɏ��J�yE_!�_%�|�z�c��̍j�_ .>��0�V�Ѭ�h6��ڋ�������������f�o/[>xZT/H��M3�=6�?V/A�
��������׀z�a��A�Qݜc�wI�� h{Ɉ�A�O���	v���d:��Dl�c�0�?Q�ڬHL޸�5[,�E���R��9њ;f��jq}H�f����K�)�twd�X��! 8�|��Q�8�|�]1:U+.b�����`ʂ���!��h�W���Y#:~S)51�ѐB�U>Q|��|l9
�}�O�V1I�ˡ�����?.Z���om7&~(ʀ�������"D?'9�@�.�\���^_�@��4��-{�%$�l�]\��Z<Y��9����sh�YF!8E�<�8a��@D�Fn��?�pw�/{hJz��lu����B{(n�v�3��!"=�)(e�����M�_熎�1l�x$<��p�z�V�痏3����1��$W��ݽݨ��KA�DH�\����J� �@��gs�jخ�|��|�az���� ���qL|�u��c�m��*�V�fنY�-lw�����k�����`�����#R��ׁ*W��"��_��!9 @]�ɭH�܀��X�q��o�?q`���Po��E�2����+n������X�<!��z�	��bf'eVͅ����<��VJi��X�#Ϡ��?����M��]��ҵ�;�oh��7q�� �>Yo�_R��3JF�(�0�S�<x�b9ʰ�JW�5 %gk(�&<�@5�u"�&�]qB� �&�n<�c�吠���J5�UN���� �i0�bgJ���r/i�b����4�X����h��ʨ9Ja#����ϥ�A
�	���!�"N��[}Le�(��Ȳ�	�C%��ʓ!�&�Y��UN�5).����ѠXϣJL��f���� ��]��m��x�Z���/�}�/@0��t
3�\�Iԙ�� �K���Px��IR�*=W��p�Y3E�.�YC������i4��l��m,M�ǺX9o�WR���n Y����CE�3���E7t�C�p�-�ͳ����u7s&X�X7�� '_�f_����@�� ��nI,�^�6m�<�Q�.�Mپw;y�Xr���=�?�I�a��-3��	 '�
m�ŭ�g�?���i�����WV^�Ÿ���E�"I��pt����&��쇜�s����>cm�	�_����U��w[�iU����+]��v��:��y��fy{��#����Dv�Q4���^�:Z'��V���3���1����~ќ>Np����+#^d�*�D�Q��v��,�)�IV��F�Q%�d���xʖ���;��Z��l��s�r>R0��O]�@�����:ʇ^S�8�O�0���k�:�_��	�r��߉�8�t��/��KP�����Y��5�Ns+�4�I�0���D��5'��	��(�ܰ�bܜ�N���Gp���m�=ǐ1�`"<g��M
ww%�"&��������.�8���vU����xZʯH}���Ƭ��;khG��_�	�b���1p����ޖ�������V�bY�Q���� �E��%'�z ���$T,��t�(�uo��>XT�3��l��bM^�,�À�����|�x��,�6�f����W'�xx�����xw#����"�
��߂�k[*3�pM�"�e�L������ݮ襘�
0w�%�T�I3?ę��u���%�.e�J`.!��;x��F��e�JE����F^7�%*fT�����L�r�HV#���0�
hve�z$�e�<VCbq��˒�B3�{��t�j}|�� >N�g�p�#�pCl�	&TCf��ى�}�k��>ҊpL�4��-���L3S"aJ�CƮ��C���R�v��:d���f|��Fv!��*e�@�d�V��*��m>�����d���h�Ͼ:e���gtC[7�y����B8�̙Y��jl�bk���k:�c�gō��h���!��6��T�zB�X����K������_�bȸ���t��)�lvi�b���n��b��M:,H���}��a{'���C��4�ϛ�e�w�.p��M���O��m�^�!l��SS�zH]J~�U�<@��B�����j-T$�/!�k��N�Ҙv"�e�xu9����,�*�Ʈ5K6~.p�ǂ�ǌ�5��˷�2#���N�Pe#�b�'PYM���ى0��d
q��{�"J�3��q������?�Ϊ���lN+�0�Z`��ذ��罡+�8�PacW�u�8:H��9u�LI�Wr}�nut�:Z��[��lk�;H�ZIF�_�
��@�k��}k���k��#�L��u�Y>��c�ZJ.��ZaH���d���]9�%��A4�ڻ��F`s$�>]l�a��Xg1����Y�\���mλ�-�՝B��ǽKb��v�!Q͹�����X�؛�����lq�#��e�La�"�#5�}T`�qf��G󨹪�y3gN�%�$�6sy0��s�`�W��MC?�%��u�|����µ�6��8�.���ҋ��>a��	��3�@����1����t�!y��8E���ͣ�_�~=��XC}�z6�g�@�$=�?�
�!B��	��w�� �sQp)�Ɋ~�U���8���ܒ�_�����I�-���9�p��S57j�.r=�2"�RM�$C���c����-vfo��f<0NoL�"p۔��MCq�VE�a�
�{!��l��1��6�d��K�5pl�I�f�k+.��|���^%:�&%
׍�Y1�A�]��1YQN��+e���^�\&���#5��b
��C�X�K�|�8������S�� �r_a%����o�>UH\�Q�A�G�-��TY�A���l��0S��>�B]l�)~W)\����0J��~� �v��0�6��&�x$K����1�Y���������t�!>������/z9��h7;	
���Y� ��W'`a�?1��u��s���$i�,ʁ�s�h��G��L�2�i({�[s��3J�kW����*E^DU`��ő)qNB�!&��F�1�)q|�6�y�28>kه@���Y�i�m�XiL��T��Y� �+���2�'��J*s��{J��s�"t�@6&$
�c����d��q�4&M�r�ƚ�b$�c㟼�0j;�_�9���=_5k�$Um�6�,,ԴRvPDi��[�3� c�8���IU���A{��=ǼHڇ��i��*��.)�S �4��Xf�Lw��P�.BoOh
�]�|AT�b��� ��:pm`�fS*J~��^�U{�;׌0#��ճF�� �����}"��;:`�40����� vF�9�.�� �b��[5 �E���wL�O������+�-�~L#0���h�B�z)��q��T�����y��y�A
"aj���=��ǒ�Ch͖��pL��`0�h*&%����-�r�M�µ!�	�_�Ѹ�e���n���/F�o ���@�wγ�qXt-�5a��v�P�#R���huE�٭O'@;��3�s�wƐ篵^I�Je|�Z�n7_���8��Y��fm2^`n�ȪF�����@���y� ��T)<�����J�A{D��nS%�>���W���/L���z�9U���G!R\6YyM�h����(��0�G�>,x��aBB�޽p��l*	?ͪ֟C�psҺ�=l�͍�/�
�]��^I0��K���İہN�(e˼�v��8�6�����!0�p��;~�����n?���J�w�y?��o������1tV�I���|
�&�bvf��{�ڹYkc��`ɣa��Dԯ#l�[xd�,gy��Q��п��C6s�@4�d�
)��c��������K,���t��)7�[�d�F6}����}����U�|\�Ɠ����(�IMͺs1�rq�p(��i;�_�-e�5Փ�F]M������8�:]Ě�ec�ۯ|Ғ�R��'��ICi�j�B#�������zo$�Rg�omf���w���g�>ڴ���2�<IQ�W��e�S*2�;!�΄%{ͪ1�zO'�N�Zv�U�r'c K�գ�0��Y57��S�v�d��8��f�U��K�q�ӆ	Lϗ�o���Z���%��[����M���o��$��u{�^����~s�Y�9�mwaH�CP�����o0: ����g/%+L�?&��}4�2],�������![�Z�!]�p%�yt�v�Kh��ʢ�=55����Ies|��i�����Z��K�����ȋ�n������__��k��-
���6��`R���I�]�O�.���%o� tj��c�z������D�0%�kt��Ʊ�N���Cz5�g8�YAu�����!�����* �"~&#`L���� 9C�5$� d��m-}���{l��!e]=\��쨗��8��C��RP�	���](�Q�S)�[��^6���U��e!���7���?/\gl��|-�m	ϐ1�(�os��-��������,CJ{s�"a+��~���]�������N\CL�`��9W�2m.泧�S,[?�Z���=Gג�� �=��7�z���c��F6[��Z��
)���z�C~K֢��Q�O�x/Lpo�?�L2T�!� C���k��Y��?8|���q��r�חC!�w>{O��0�3Y���y�y�,k-*��+� l�v�[�c$H �e����>��^Ww�3=g/�-G(I�͞�_��'�}��S����;����]��N��:��w�e�d��M9S���Y�f�d���o�9?!\� 8��>:z���(s�/����Kq����i�l?qlu�#6 �^�77#�`��k���,E���^D	��Zn��"�}�n⁹�^�����Y�_]QKk��G#����²0�W|���l�;�p�H�#��H��nv+*5�7��l'���;	gP��b��[0T�b���粻�X���'�2�%���i�lbٖZ��q#X�������5�D��*1�����#��9ޠ����4]�>�g���ذprx�iR���V:-R��?�B���	�s�;�_?ɴ�����Ӷp����~2P$¸PlPsL�����Ձ�q��Q�)��Q�;�v�� $5��7j܃�������T���N�vN3AA��� ���	�6_OK+?Q�}Ҙ���[�!O�L�2?C�S�M���wӑ�)Y��S3/m�R�=�c�Tr�مmT{x1BV� X����{9�#ٽ�~W� <ż�dK�ЌfnOF�M�$a�59���O�+n��1o������z�LE����;s�h�G*kq�EEw"�?������_�q8�?)�B��G
���J�j�g�qZ#j�7��t�?����"w��"��!�)�]Q����u��X�(�Ac�\�'~�7�e��C#�X���`�����u�a�B���,v?����k!�?��J�v+�v�B�t0Gg,�ʺ ��VN��)q�@X�%�e2�&A�#̊�q�����K��I~9 aV�r_laB�4���*U�؈�6HIm���<�)��(����>�L���o��v���0�I��>�]Bq2� ����YH�����!�i�*���t�)q��ܛ{����9����]SI��y]����oF4�ݹ	��*�ڹ�T�_3Z�<I'r���lCh�%�^���Uؓ"���㒟�jm�{��!�>&�2��<�߷���uC�6}^�7�4���|r���%V ���털��ܦ,�<^��b9�0�(�#���'[��e�l+��Ը�y���j0�t��v��L%�e������N��(�|j[��@i�l��ZA�y����~i݉z.������pr&��p^�:���]�@�-���t��Ʉ���xU���Q SQcQ�к���_AVcL�+�1�iJ���@3j�#�����@
S{DQU?7�!r=qGɭ�P��Ȱ�q�-��RN�R3�6�s�z�����b�v�|�~bi�]�&����f�F�����a�31�w�X��y�r�ar@Q¾�|�C�!E�9�ج�\r��%�t�v�<wb`��M����4a�0��7M��-'�8f9�)�Z@�}���$�Sx[�cD�A�C�����U�����5�L�X��W|<����J�Q����������?{��d1A��$A*ݺ��چ9���ZTS��pB�����L��ʢ,?P�鸤��e뽚� q)�F2�s�o��m��Sԟ�7LP�����߂5a`OKH"����c%�'a�|jmU�s��TqN ;�Vw�3�Ps@���d�%�u���W�Z�?�H�	Ńui�n42�	��E�ڟ
`�7�.���Y̐�,ѓ;�s^L@���f��'c�f!�����R���ډ�!j�N=��@ڵ�gMX�گ̋���CӀY��I�+75��s0���&\
/�u��K0}� t�Җ�_��.��;'@����t�J�6���JVB������e�V�X����M�
�/y~P�79���Uh��,��h�)�>c��8Jk?�hb�� ��6���6�3kL}�Q|G��(�7i��\����r�n9����~��$ID�5/XLuずQ�M�A�ta�!̭�H�Q�!�5�	'�)�<E�
]K��O>!W�c��y���N��	�
��vӮ"�j�.��x�y���y�u�*V#��Ґ�$1"����!׸O#}M��S?��V�Yd���V0����,(ߨ;p�rp4��+�����`Qc\�{|[-� n��MI1��Cr�$x���������@r3��ઌ����ZQ�o�y[E�=ҡ�"U)S�R\�<�u��+r@��1A\�y(�de���{J��S����x$�2b��|��7 U�M�/���b�����yO����Ԩ�W\t��^�%�r\�Te|����N>�ZxI�|e��%��\���*e⧯�$Q�yfH ����6�J.��������{u�C�-�E�8��#;�Z��ci>��b`h�I)�e�7�E龧j�����k�~Gl�w������=�P��Ԭ�Qg�����]����$��bߝG�9��v�����.�MQ^(p���T�B�'�M�C7ig� ��rS�[Q���(��aHZ~�X�(g+ǖ����Y��#�Ƃ��[T�9�% �OY	!�5Տ�7�����l"��������5�����#��'F��.��/�UGr�`��l�٫:$h�q,*W1�9/���D,��FLH����n~\*�˟�m���ܧ�����lS⇳0�}�m �R�f�Bㅫ���e��Luc��]�1j�]�H���²q�N��rn�y��|�]a��n�oKU�'��kQ�;ͷ V��VJX����L�`�d��~?�X$!~8�ƈ���%���tDxS�HʔT?B8�Y�����YO볶O��[{;U��ץ�}Q�J����VH&�������f'v��(f�q��.I���g�/�I�"�]�ѱ��0l�g�0;���nV�⹁<G�c��y%9��#`��Y@���N�n���3˨������.���Ԅ�߾V��}A�z��*�D�iؾeAA�p����%bɚ��Q��{�-5����i�1���r�$�vs�K*��k&	���D8���]$ ����y ��"p%n�W5`N��%ר�qp�όL{K,���K�(�Fl����G����$>-�;��L1�{�����+�2��Q;��	�E�d���	���?���O�:����E���O���+����&J���"��C��Ps�����*$*��̽S w��"��D�E��?W��OJ�+)ٶ%�eq	�T���_o��V�HaՆO�=��:c{0��SD��ʩ��8��ޡ�"8M\/�l')~��Q/C��Q���4�Jj�����8�_�����EKS�K2���2I_M���mT���5�$����H�
{@��}Σ߉Y���?���g�����n��aU�1��X��]$"�`:fci�+n� I� �hf��;TF�|?�@��.��7�H�h�M-S��������A�˘��)��FOB���6jl�x���0lm���Hyx�\7�2��t@��{�4{V�S��ʼ��
��]�`c㍬�����!��
���R�w�8��{��v)�0�#��:����T�n�n�/2w�kl�rAǠܟ��Ku-ǯ%���-.N�U-V'h��UΩ��YDw�EU� /\��Qc5��3��r�ʚM���B\�-��i�Sa�n�P�����Ax1�gƁ ʉ*y�o����x�q��vj-�uRo�
�*��R�g�:�J�-SR��&��f�w�r,�ԣ^Y���B����8F�c��#�'�O�A�������p�d�%F�U�W HI8��o�j�9�^�ɸ��eRnޏ�B�M��Ycw=5؜��ף`!�>#Ӓ.2�#GD(�6oiT���i_��)ZJT�PDa	��������MɬE�C:�BqЩ���P[�������+�Z���rDLLB�D]fܼz3����-��N>��Lx�g���bP�M]i��i/"El�RM��ٰ� ����$^�#S��Cé�����S���O���``\?���]ɻ�ó����x��󛧬�;r�H�l��	z�d���H0�и�^��=L�q�+k�t��'�D��|�EZk�`�0N�7*�6��%KJxx�ae��8�Ѱ��E�v�F|,uso[٠;8�B�=�s'��S��&ן��F�l��7P�݆���ش��a��8�ŕ^�m7.�8���"����r�썃]�.ϥuȺ8��Zĳ?�T�������G��[�vJ&	x��6=o������˅Ì���t�X�<�F����U�3��C�]j!������/\�3ԟE�N��Lҷ��-�o8���q�)П�{�E��E�20��R�K7_v]:��iAd#E���#{�-7M�!� �&�j������)#ֆ]���;R��C���}`�)�t�f����u҇|��!�v�6L�xY�@�ܷ��x���FN�Y�uE[u'��-�y�L<�z�4D-�ˆ�t֋�u��E Rz-$��u&'�+���k��#{��pT�&}!C��>�������r��('���
f��)L�Dwi��WayS��Hp�mBĜ�	�$����
�le�L0 J����N�.�4�_
wR|]�a-X�L��
++��(�د^ɍ]���,	�~� �h�#��Iw�
q��V�W�"	��B���~m�T�<�*�ۦ�W�I����d���料K /*n�&�z��Gb���QbdcAy��Q�!D)΂��#�5�O�c�&٥,]��;T��ݐc�����. q͂���X��M��@�pr��e7)$���p/J`c�MڇA,_�&k~Ք��g�q[�+eT�ޠ~~[��9w�t�����s�!g�U�����*��z�t��D�l,B-t��|*M�����M/=wiØ1t�N�6�835�Cb��Z�*(�p�`38�Y��]�̮#`c�9F��4?�#��e���,R��]zSb��b�J�� �]	�J�°�o�N�$V���]_��Y�C{�:�����J�t|�W.�	�X�������[�b�MA�o¶�W��V��,`���ojK^?�'*�MH;��� i܅QU�"�+X��'��C�ţ�E��:������Ư�jV+��4�%~āОٴ/���m�&�ߙKMT�)?����&�-�H��4�;�=�6
fL[4)�����h���{��Lw��$�M\WPՀyb& >7�����H�
uD��ٹ�S�O�2��Wtm�#�	�}'wsj���q㛮s�˺ơ"�S%�P�G�쪁H��q�;e�?���N�.)J����v磉����J7�H��M����n�����$�����T�wu�MN���G_	o�[б�6cۋ���<��5�1� 6��}2�����y�� ��Jm�P/�T:�/XAҌ`Jr!����w	����yz���:��M�.��~]aLb��hh�ϒg�!�ցg	#_������~W�4l����fM/��H���K�h�IEg��Ҽ��F`%��\��S�w�PȂ	��y9�1t��;��@6d.�A<	��m��8]is~������E�^��Zh�X�P��=R����l);hn/~��/��q�G"�G	���6{ �{z�w�$���hȾ�t�G�	Ԃl=�!�N/%����祇�ߎ]�K됎i��Xb<�V��-�'N]��z)K��U�j�>���$�q�֑�f`�q�eRW�֬־d�U�As�'�E��-O�D͏*�?BEm��z-@���3 ��mR���z�E�V-�_���� <�k+T�A�;ܖ�H��[�bI>���@M���f��Bz��Mh�������+ I�,��g t�1G�p�+���)�n�J*���%��E�+2e+4z��1Ȳ�����J�(#��j��g�؊�(�������	cĮ��@@�� �5�U<�������`�nӣB7
1O+
˵E4���l�iD�^�.RQ���g��+�G:bז�і�B�.!�w"�i�M�e��B#����vׂ��f��P<v��ܕi��˝~f�y�鴒FD��ˇ+��E��N������
����KV��&����a$�rQ,f|��-�����"�9��Țё��j�F��7J�g�&xH�i���\�a WK��8�&�t�t�g7N ���m>;��L�#�_�N��oz-j�n�Wh)��1�ӯ���yp<w�c��)�|��������F!Wp1ϱFȣ	h���9�F�����_��!�W<I�?1�V���ƼS�`�QRy��d�ɾ�G�M��p�jR#i�jq����t�<��g�����N#�j){` ��~�W��wQ�ch#2.�e��uEpQx�u��QC&�u�X�����-bS���zػ/i�[��֋=��4�<-J����V��#���W�k�(ǸC\K����'=���dR��xאz�����S9P.��d��	����<�I����Dc֐�\n����̒ǳ
�6������7� X�9�(c�0�~.��� ��7���Nv'�8��t���͊=U��<8LE՟��MnϤ#�Xn���m���[4fb���o�_��v�A��mÍ���Xod����R��%@������;�B>{����؃P�B���i���zO��ǖ���w'k�;��o���7�4��;E�DG_��l_l�1}[�Ǧ��`%�\oI_CЎҡN�^��:n�4@�v��O�{-��E)(�|2m?UR`NzD�t;��� j���Ϻ���ߕ��'��e�!>y�	�s�9�Xy4P"FaALQ�y����x۞�P3��@A�E�(�A WQ����X�=w���w�����s^#�c���f�C��^��m	#y�z��� ��?���cd�bOC9*|Z�ƕi�8�dI꺳Ѝ��Af�.û(C�`c�4����:J{��m{��5���fM��m��{��2�Lx
?QB�?O�h�. I<�H��-�4uIj��^���鬣�B��r{�l���/zqc�7���ѼF�ivp4.TY]�zp�P�US�	�OY'��"�뒰��ݵ	�H��ǡ�^���e�M��y�
n�\⇓yd�>mݳ����]?���	����gF9� ���8zk���h#���2ot�"쯩ێ�αZ����� 	\�`�H(����J�'5t?o$�|�"Ge�xi@�U:*�
���W�!7�K@�_\�1\��� �J{r�D�i��_�4�`�V��͊�VqdZ�o"~�V%�����D]��f?y���m�"�J�rB�!lt�l�qy�	~��Ǌ:03"�?�s�ŕhՄ��98a��줸.��o�_������i��N@���:�ݐ�Z�8��#��1s�����:p��:��H:�{�77���R:븂��~~kJ_���<�ڑ/�G�<Gf�[G�����I�)0N��K�D�ļLR�U���&K��W���Z�|=ѣ�ˏ�9�I�1�]���������69������T$d,��B��c�ʛ�N���9�@�RO����G\C�bA�"�$A�����Sɀ��y3y,I}�U�"	�K�GR�r�va?$� ��l�7��Zuz�0&��[Bã^@X�|3�����ܴ�y��ɞ��VYr&����	_�]�8�INM��݈|�ݿ�p�fl�������Z<�X��N6z�ԭ[8��|}�� �'/(:�/��}�)�脡��݄���E+�{��GV�� ���٩źZ(��c�����^�o�<��GJ�B���Q�U�B�/�Dd��F�zY��9����L�GǿA���U̓ooDU:~[�4EbW�m�� vE�1v�q͉�r��uڀ�邇�dYSq�2 ]��i(jh�'��4yL����3'̙�F�Y��]��O��PM,Vz�9���/wb�����=򜨹���I�zBJ��V��Kȴ	�*��}��ݮ�j}�6���І3P�������}&�y�Ԟְ��V�zrMrS��ژ��I����V������s7w�'i"s�A����Q��]Z�����ö,ei���������U�Z��kAg����d9����+�(�*o���lJ8y�!�S�L��G*�ί�%W0���D�����$��v43D�GWz4d���';���6���`ɚ��9�fC�Kl�̒�D�l1+Ƃ���<�XY�sL����n���EN�tYP�mQ:vwg���˙y�܋d/�͓b����T�f:���6�"f΋�Ü�R�/na�> ��QK����rJ��Wo5�+��MF$k)
w�-����ԭ��	�D4�y�5O/,�U�O�F9��8���2_g T\6h4:D|��0[�Ψ��zO��o�է������*.ZLX|z��ɯz�H���h��	�O{j*�Y�6iɒ����;���\��5�O��CĪ�>c�;��]B��A�3�H��������J<�ݽ�,Î'��M����X�-՞�l�~�J`Qɣ,�(�B��^�S���EZ[���ѽ���<@9T뮁�	* ��Ь��Wĥ�h��������7ȧ.����R�̜ߖ1�Y�#3�B		�#Y�U��O�w*��?@� ��M�~���:<���������ܭr/���Ri!H@;ɝ@��AV�g3�m�"M.70C�R�"7k�D����hP�hvSqj� f���;O}�g&N,�7m���;x4٠ũ�pfi�wFm�819@�^��Ḍ��'�ÿ9H@�*���>y����Z�O�`���w,����M�5mǔ�i�3ɰ5O��w�Ж���ٮ7	�Gy\�mpw]|�`�@�\+�,�`�q�hi�4΢&��]����,'}�Vb�o� � �.%���^�:�S�:�����17����8�P;�G�w�Ĕ�&�'y!T��������Y��S#�'WeO�\��]�o*��Np�2���%��� Xu�� � $eE\B�L�%��}��'����lbI���_��.9���'ig�Z��=M/�4��l(h��Pڲ�Df��1�������?�����#t.y
��������d�ܶA#ɨ��@iaC�_qE|���Ք&uv�[�=8�8�����?dYπc�#�u�6�D@e}�J�_9۵�;H�����i��ϱx\Hb��GЧ��@J��cċcq�ε6�لmd�6�x��@�
^�X��v<:������I���^��?R�����Ō	ޜ�}�����]�J���|���w��C4�%I=⻃�y�A\	��)�+HwD �#I��-�z�K��s�[LЕ4���[���O���?o��z�_�7��������˰&W�6��w%�ԧ6"�����b�<�׊l`I���Qx��4�|v��]�]�7D�:RXT���d^}�T��}Ҍ1ԗ���� [�o�G��VY4ZH��xujA5�|A���Ny���h)�p�	e�� �wb��e�WP��]�k�p]r��JG�P�'�$�OT&kNYNT�iC�< 3Y�7�ґİf� >\�܆<�(��乗��wn��-��W_��ګ����Y]���8(�~@�)Up�����$���%{��vnN07���K��u�3Ē��4o��X�w2������]7�P�[��L���R9��S>�Ĺ�o�ѹ�IS`�<��Z��z�¯+�z�4E����x'�Q:p*�8��kDa0*��-�vd���u?"�]Ev,��wꅼ�Ѷԏ�̅V�gL�  H��gu���F��g�r����8�I�B��,�qQ�ȶ/�?:�-�B�I�ټ�[(ʓ/'�{/%���[OTh�=�5���S����F�c` ��i�^�f��K�V���/����y�t79K�������p�Y��ƌi�C�� ��1Vµ\�%�;�5ܐ����`��7Lf��k���N���c"&�r�*�WN�����c�zx�Ơ�(��&	�,�@��v��<p�US>.Ĩy%�r�����-Kk�_����H�O(pP;����r��lu��x:?+�*0Zr���~~i���Vd����<Ec�.��?��@V�(�|�&���H���[��_�7$�n�@����}�G�0G)6�Il�:��m��$ ��g�c���������T����{
j�]�V�I9��\���w�gne昸c�Co���,�����oJ2��b�4�p��$�˙�k�j�+�U?31�n�ᾙQF�20�vcbH��2��8�V�K��;�R�
�u��`Z=��Q.���� u{p�[:4F�R�L��A��B@�'�����b(|����5s�l:����9�|�5<u�m�tH��ܢ��>a3eX��� ��)fa@���N��i�mN,��O.a">��ӌ��\Vw�,��U���Xה���J1<h�Rf��U����$����(�Ot�Tܱu��_��f�&��d�� lI��ܕ=f��D����!��4p�����Cxפ}w�����{RDǠV���ITXÓ�	 I/e��vk�v�c�mr
{��V��yu�,BS���b�y8��N���>�Ԛt�����x�,9$�����Ǳ�s(ܸp�]ͣ"����X�,�- ַ�qP')&�e)`Ϋe4���^�f�!�7�!7����]���^H�A�ONYi)���N��bM������`s�%���QSk�HK����,A��e�l>�ʲDF�+��ļ���ǫ%�4�T?�{�2U�A��������v4h��$��_kP�-=����e�r���������feȲ�m�v��i�=j����9���H4V7�yi��č$��}���"�k����Z��VǢ�h� G(�2Ȉ%̈�t/�z�,�3�C5��U`+f�g�@T(Gf�q��$N��3�ġo��zQ�����5Q!�!�g��~����D���(i�TF:���[��RC�CS�S���X;�l}��nxKx�$���?:Gg�w�i��Bx�� &�6����vd���-�!K�*��@{a���x��,��9��U��iGx�v�]ɾ�ѹ&�I��Whg�.nZ�V�`�<�Zr�145��Yz�{�\�ĳQ�OS��~�P*��zuY}Q��,��;�f٪L
K�zK�����؄$�tS3�Hn�����EIܠګ��܎���UQ�t<v��|Cl	��cP7�=j��Ѡ�=]�b)���RQ�&VzL�~ȀV_}i7�����1G?װ��!�!^���)�a�L	�2�H�E��	]�����>"��^�r�_�2>ٝuV��d��lT���-��xB��M�?����b��V�v��9��׻Ԑ�Y/.kE��%��z�hݢ?l-��NP�_-M�B��1h�ɥ�~���6&����-�~�1=.(���-�`�����uh�\!��|���
Ϝ��2(/	"���C`���c��N�c"h�$�7� �`*�c(�;�$H~r�k��7$�S)6�HZ����TKƖ��
C��Np(V�fh����B���qQ�hp-��|[��T%`!vN�GX�ki�o��ҁ��u��i5�ԉ���,�\���`����9W�����o�X�m�#ë������M���M��{���V8s��u��@,�jwI>
o隡��{Xe�a����w��U}f*��[d��g��f���e��h�)�;���arI��z�M�_#2=����5�xx�K����dsa���L`�y��P�JC,Nb��N����yizg�"S�m~�i~�fV�D1� I�_ �}�c��d�lv*�*��0CA�Lc/���= e�8�Q�zp�E�s���}(�*��0��
�X꽖�O� }`iu��H�Y���
C�9��R9͌�d,�H*d^I$��q���7	H�'8�1w�A��I�����8��X|�U�]�Ԋ�.�;��Oy�D�י��e��j���R!���Þ�LGJ��7ա�"a�5�c:*�K�í&�} 6�J������7&(�=f�Ι�����xډ���L?���dwA$��Uih�;r�@�~j�䊃�mc�B��ȿ �K-
:$�蟡X
5�w�U���p�=�I�.�+/I9�{�J^�(�=��֋�܉����2^ɷ
S�?�`�u��[]"�9h��#y��\�Հ��bA�zW��t�9B����y�o�%_&0��Z�(�m��_��7�T��'}D�AL�w&��n�d&�1��	��kE|�"z�1$����IW�L��zk��]ٿG~8�ƪL,BZ�=g4�M!��MA�-��Fi�O#�;��*�8N��C�֤n`E]��hJ�<7�V�1�T��.#R�Q�0�f߫�%4���0�b�QgE�(��S�i)�g��^c�%p�=�ăE��xVNLR�A��7�{���D�n��hc6zX)7�Sҕ���F<ʟ�FR���<�������QR]�T�w"�VA;�Heo#e� ��@�q������,e�Y���(�J���i����+�5+g�W�93�k�������74��~� |d��6�[�;4z���>��� OmR��E}�5���jp&��U՞��U�s���2��E�~4�tM23 ~���G�CD�$��I�E��D��5~��A�v�4%{�ꥴ�>��<֪;��V�5/G�5��7��_F�z5�t��"r�QF�E���Xq�ntg^�Ϊ�Ec9��=b��._���$;\dut/=%P�쥅���Q��J/w炙��R! ������2�(q���Mu��[�Q!���aI��]z������E Oq�p�h�T�v����n��<Jw͠9>?y���'KxU1��$	�5e�������"�W�l�e����W��nZQ�A��� p�y�jTθ��v����+�ȍ�y�U��kZ�3���kRq��i��J؎H�4͂�C�~��z�.cn,��O�ġV�2Qi/��(�l�X��L!M�T;"�y�AGw~��z����A*�����P�j�s�>6�C��G�&���{��>rxΘc��"���� W�ֈH��v'hF�Y/�X�h��v��<o�!��@]jhN���3���ZA��s>��1�&y<�hm�=���>zf~1��:/&c;���Tg
��RR���2xB[9T���M�帲a��ICL��L����u���-�� QUO�����Tc��!����O���`+��	>����K[f�P�䅎w��$�V��}��{��a�#�"G]l'J�s*iP��ԟ�q��f`:���*7��#"����߯��[�����U��_{� ��=~�Z-;�%��8���� �;��_"����`8���/]��(%�3���g��%���>�٠��T�����F�1���D/�'J���ͳ�v+)����Ÿ��
څ��T�#l\tO]Yt����p2�x��'z܅j�\�SՉ?#wK\[LmPzh@�o��0.� gi����թ��)v���Ζc�t&������!���i,~�H��LF�i���(Vv��3����4Z�آ";(�@���o�R���������í�Q�p6��K3��&�\W�u����_��$p���������q��A�]��3=纰��v�.���z����(�A,���֒b�R���ޏ0��$>�ߛ<���[�}�tz��5��V�M!߽'���(D6u�S(�k�9��u	����`�<��ơRqXg��vs��Җ}7��^ؾ.`����8�Q�����+�H��ʿ��1���.~��T����5$��r��eO]z�3��$ a&�	���&la��qL`o�Q�j)��R=�\.i?�̭b���L�~K��el*N�^3�n�}��Ro��γ�e�Y��$���7�#K��em*Gݬ�ýa�#d�(���iV��@%V>�&`���z�	�B{G)n�V�����!ǵ9�A��&�E�������Ki�i���P�����1@r�/�);�	�8҇z/Va�� m0�{�O�
���a&�*�ǵ��Q��+|(ɩWFçlx�Oq?W ���QS�d�Lɧc"��pYwȠ��(��8E�GdH�nL:|X� @^��"0�
�y�(d:vC���2c7bt���s��:(��z�*uQ���	��+M��Â� ?�,�Dz-@�OѾ�.O}q�i0�G�����g.�\�Ӌ=e���]����	�ŔXǱ��El�&��bW����P�U��P�m��ʥ�t����������z�k����JE2�%R�M�*@9zb}B�21i1�ڵ�J�A�_�y��&�E��J���`r��MZ��>"⤍ �ƕ{���.��@���~[����o%TF2��wS㡟�����),�6���58���x��/���cƶA3�I��H�ro#fw
[��G��~WS�����6ְ��;��96���3k�g΂U�bй�P���&�>I߼Z��f�fK/��r\a�<U<��=�f�[x�,�p����l�_�fG$������P؊S7�/�<�ԥ F��b�Wx�s��xY_�h:��n��fcvH䷒͎N� ������Kd�Z_���ߓ8��5'�d��~sG���ɵ��4����׺@�:�*�NN��7�ǅ�b�K5�_�� ��.?�9�_\]s�����`�[�<�Eg<ڱ�P.-y�R��A7J��x�/��<t�\dA�n'��t��L|XY3���$^q�i�dz���XXz�t��!�=��h���K��Oz�P��	ު�%��6�Ɲ���窢S��0/ڃ�3Q�b���X�i���]�F,w$���(Rv'`���BYlWO���ϵl��t�Qɺ�3���3���yP�����R%U2�[���yNeDY��7�r�3���4@��1p�HQ��X��[41t����ݻ�P1��ܰ���U
r�х������1o7�#���Qd���� ��Rx�5�StW��y�'(��0���@A��a>�2`�i�XO������
w�M�S0S���aX����vm@�������ى�AT���x��E׌���`�Ky5M]p�yg�!(u��5���{ż�p���B�B:���ԇ*'\�wj+�,�fby���
� �#����5����X��f��5#��!~��^�H7zw�]��.b�[j(�і��D�ȣ�C���L*�퍹� -�g�-��[,���<��1*��۠�;L��Eg^O��F��Y�����&�sKd2ۅT��vT���9��-� [�N�R{r3���u�r�PL�Fd2_����`�"��������\ �H���.*�*��
��|�M�Za����Gx�G8$aWq��\�|D����e���~r�9��ou(�<�Pj��Jc��<��tI?�=T���vY�cI�Ϥ7&>1	�[sܚ6�*�B�(2$yl%ı��z� ���p@����Sʺ���1��IS���E�.�+ Mw��[w����g��5�����n�Y�K� 7ܤ'L�~�>"��ʿ}Q�Ο�O� ����GbB�J���(��T�	E����㦼&I�x5C\wZ)�F+~��g^Htm���3�<?�F�G
�R����ߺA���kS�����H�\��#h�t���7�l�*}�+j��Z�҇��)�(�l�P�xj7�����ݙ㯈�X�dW���Ӹ�U'�)�(�U�v�4���wR;��/��:ױl4���<{���l�g�1�fiC���:�1a\����ݳ0"+oQ��z_.x�I2��HCڢ�+�#�*�3���e�� j�LBݛF�ϰݝ
�R�8�����x'3�����D��?g���1���V���R��Ț:�'у�����q��:PY����Ͼ,Pa�������~�� ��D��gy=��^�&��.�䕁0�����*4pP�.iR�R�"�u'J����}�}F��:�㲴s�5�|��aϱ�_'�A�R˅�V]&��\e���˶�׮3�5e�ԓ�#�:cm��%���ᓹ��5�,}��xVM�"R�zR��e��dW��V&v��tY���ISy�*IYY8�����?�~_�|�ʦ�n���I�X/}h6*�q0�3�2�-�P����CJ+0@ J}��x�rO�q�{p��cw%+�K�{�GW�2g4.�r5��Y\�{��IX�_����o����e;TH��U�hʧe�Y��Z�\��R�F<Ql_ �2t8�KwGa�H=L���`p���K���Κ#Bɇ-9�P$�0����RZ�����#t�c�����C��/�C}��i�F���J�e��7�ۀ4i,�u��s��e�r-�G�NnUA��j|`� �R��Mo����;�����sa�ʇ�n�?��J�_4:gXv`�	�=�Wյ��N�iЬ�=��h��I	eɝ!�sc����~�3��HR�*��Sc� ]#�D���>��u\Y��YF�Ꮔom3���U�H���~Xt��k*+iMuF=�h˟6�-2��"B�=��tK2p=����z!���W-��Ns������y)��)�nB�H��l{T���Ru�64L���u�,b�3:Z�s���d�+lZ�u�������h��̼���$��~� �O(�iͅP	]Q)��j�o'i«�Y����m�p��z��;�`��c�A�S8q�̠�$�$��@"�מ���$r�2�~N���<�M��rC\�3�T��^�.���FC�*fJ�x��ˉQ/�������J�/��컫�/���P=\gL휌�$�qZ�M���� �SX1�.�!���k����w��ɪ`=�d������A�G}4	�&h��R&�Z�}������b���\~ �!�Se�����"����WJ,n����M���MkՐ0l�S�d�옑$�5�v���N�u���Q//V�`i�aev�W�B�6�H��wS��Q�V�Ǹ^��s�_L,��d�Y���}�օ*P�\�]5��:jMI؛h|툓O���}SCS��ې���M��az�UF1�
hݷ�`$�l�(R�ֺ�-,�8kl����,��u���RԺ�OZҜvm (����P@�S�~Y���`�$w�t-|����p���yQ�4b��_6�0�� ��kMQ�lA�|��h�Dy� ͙R}]�{��:��N ǲ�J�����ڑ��,�-)�_q�wY�G7h>�� �G.��;߹��ջ�k�!i���q�1�^��ͻ�b@u���\�mT��W�@&��y{Ec���U��߁Y��>>R!��\FG���H�}�0�
"�	n%H6�AV��S���tg�L�:�=�O�Á�%7�_�-����(:��;��������2�]�˦�+����X��=9��!d���S���젌gc��ΊZF-Wp��xT��EZ-���������!�lsv3&p�'�q[zJ-�Y+*~�jFM��S���'����?�Ƭ�O�/X�t���hڒ�e�DQ	��3o��n'���O�`U�	������VY��K�5�c}��{K6�&�U}�`c��N�XB����^�[���0YL}�=���8W���SKr͈9vi�����ʣF���'"q5U߰M�Q����Ub���:�q�Dj�M�j��a���As�*�*`R�[X��҈�	���{f3O�%;��5�� d��ү�L��hP����'�
�l��'#.z��3{��Vk�
_��!������b��.����#����yͶ�å�o������*�%(���o��U;����B��C�P��� ��HF��z�3��{L�XM��P���1i������.��/nL��Ⱥ7�K�nע��N��k0�P�i�>G5���Mtj������aTs{�-�xJ䯘�.e	I�0����ݚh����vA?E�AJ���h&��VJ$�������z�g�	�c.!��,�O3�$��9ܦ�V-�}gޟ�JR�:�ф��iRC�)��8�n��C��
�O�Ce�	�;�K�����xOϧs��PA�&���3�.`�%'`%�y����Q[b0Y��4�����܈��W�U+�2f	XF�>l=7�lܚ2UV�W��I���^0�{e|��p_��.
&��ξ
���V�m}���M�75���.;�\x��5o��7i熞Ǽ���8�Q��M�]�*!x6\JXB3b[}���w�U���cO�(D��n���7�8��h��dr���G ��\�Crm���z��%3�/(w8��(?
��j�+�d"B1Ҫc+�
F���>����".�1��d�L���F�I���}�F؋��*/���y?�z����h�M@k��x|�	\�L�-��UƄ���(8�-��O�yL�6���[�=�`�x�sO.8����i�24� ��d��Q]{j��y��Z�P�샣F����ک��,.��+Ar(9ޭ�)��D�1��o,68��4/Zb��(^�FU��Nr~&���cN�%]�w�'�K�u��k�����Y����UF�j;[`�T�b2��,�N��tl��%d��6ȑ��32�V���yژڜW��������b�����9AD�v�+J�s�8�hO� ?����50�������{��
̸^���У��T ]хP$4+{�S�=#�RM��xM_߳�QH�yt~�
Ɓ�BShZf�MV~v�G�e[].@R�%�p�{b����gwp�0E*��=��2�%ΆG�>O��v�?9m��WC��/���)T�Ŀh	�gQ�����m�������0Tҳ��(�j��1g�O�{T��M��hFir�,��.@u)����/&�+�0�e-�R�ij/_�_�A�dE�B��PT�E���^���%��1�/W;��9����k@�D�T�m�OX+���O��ۮ�,f '�F\��+"��W�ܯX�t���F5��[�kah�j��aX��.|=�p ��`Q�0�3�Aĳ�k��n��ń�vX�*��Q|/�י"�r�o��9��2SKio3d	�6<�۞SV�d&�6A7���ֹ���7�L�Mq�����j�9�D,`~�7�n2
u�}��\�g��o]�dV��uĝ���*�I�uk��Q,���"Hw��Ѥ(\wX�)����'��䘆x�`3)��ߟ���/.��L�ecm�~ S�}*s$XfXH�H!eh�d��kv c�L�?z[e�g�_��괊3�����<��#  ǃ� |T_��]
?�����#6v�M�n(!��>Q,��& X��g`�%!������,N;�gPEV�b/�zZ�k�`m��}�!���v���]<rmz����\@z�ڏ�`Ʃ2�Z�U��F�4"�_�7F��O��I�b��pR�s�DƎ8�9χ�[�?��5{kxW�C���B��pL���$9IQ���nx�;���7|xB�*��q�4�Y�y�7V�d�m��9l`M��4A�O}&x���O&��fi�b��,hF������oU�� l�hש��Ƹxi�]��A=�N���)@\X�
����m��R��@FՈ����%nkXC���e�PG7����1X�Q;ٰ^�Sf=PN�����VJ�3�o��[iU$0��9�S|��L�m��c�jr�H���g'�����<��lezH_�TQ�ȡK\�Ŵ�J�t�f�VQu!���s�j�ܖ�Z �|��-�'y�9�)�I|؆��N��I+��5�®!���g2�8����0��� �?��.�c�A��,����J��y���ɶ�s��7�'1��3ao��������dcPK_~2�&�Es|�]��0��BR㟝�'���v($E
���fj�}@6�Ռ�dL������r� ��#�Ĕ�|eP�w��S�nPBy������T�Sk��R�--)b��8�� '8����>�7��Z���K/�� @&�v�8���,w`F����㔀S�fe��I�.DuQg|�Yt�|�J��Wč:���}>�VK���	h%�d�����PV`J��b+�x��OּFXz�Ô�o�w���Jd�<?;{=�r3`$wV�޷&�����A��uS��i<�t�x��fq2�Z�聠�x�a����ğ���g��P�+����ӿ��TlD��_�-$�zz�u�����	�="��]0�O��O��c�w,�c�;7f� _A���l�?�۠�����P�a �F�޴� 8�ѽ7; �a�4����1�B�Ǹ>��дD>�U��׵�>�[����ev*�J�h�Ꮌ�l*R�t�����u���o��dK�V(yvn=������<�+v���޻.Ѐ���>'O��(��hg���\�S��(,�a�b	SQ[�
ToJ�Ɵlf�n��5�ɛ�>+7�݂[�?��<���js�Ve?WD����-Æ:��7Z���M��B�M�L'Fcq�D-坝%*��M�Q����=��K#���0.���@��Nײ�&�K9͊��A�|>�eqH�%24�8'�)��	Q��B/�KjO ��$��T8!��+�+�%5��T|Z����hB�?�5�Ceۍ���3EhBH)F�_	5��ۆn8[W��)4������A!<7��T΍O�z��� ��2�U��M?��M,	�^=xn�5��Ӕ�����0J�	�3���L��o���m݌���:�
�6Mk9����e'�I��^]��L���k��%4�L� �j��τ8��3��C��qe[���kN�_JqOy�۫�} ��,&�Nb�X!�'k�0?�i������K��1]��?�V�ߴ�}�ϧ�v�)9SKl�1#��߾��lb�o�^��sүZk�-�x
mr���XQ(YR�G�'�<�Άߟ��y�8���wrٌ����򽐳�����b'�)]mm}�"f�G/���ǁ����ʈE�r5��h���ɋ ���%�z����E+�h<6bǏ�X�bC�&��e�mqrX�xb��Q�5u�F�����w�c��#�ćmb���qc��|�:�(�q�#���P���XXׂ�潣.qJG==�B6���p �i�L:@�Ci���XO|N!dLè^'a��q�ӎ�-}D�F��v�92cL���M� ��{����q��ɦ`I�����[��{	0�@�-�1� �T�eF�[H��E��d����b;��xۤm�}�Q���Y�U��p�A6�&IT-T�Iʩ^��+�uF6�G�x.���C΄��-����.����A��0:+<S�^0_����>�d�s~���<�U_~��Y����,��P��Ș2KWc��Uxl�o�N�EN!���oP�����w����_mؾ��*�����C�&>�l�wZ���9��2�+��tE]� 4)�@�<�pDg9{�
W�X�\c����?��V�Έ���5O?�l�/����yi �k
�£���w�ET	x��ׇ��*3/�U���H�N�z5ca_�??	#M���3%����u��+#�v�� �x񃌉�ĂhyUBٌ�涁`A±�
�U�N�ӑY2�h�T;F�*E*�?TLQ������ؐ3��8�a����K0J����3� ��j$�����Z-����c[q �X$]B���'���Z�.W���)�Jb��+-�Dܚ��.��4�I�v�'�����ȱ.Rs����b2�: ��X�H�������)���AM�T�1��0G���&�'·K�r˅{�dn�h
B �Sa�������1��\4��ˡ�Q�I|��3�R��j)1�1u�W���'p.�r��BH�P�XU���TT/����S?V��^z��PܼW&�E�r$F�r�,e�%^��MJd�R]Uf���Ŗ�B��Ƃ�3�;[�W.��U���<�X�<�ڧ6\j�_�T��Eq M�B}h���0��^���<6k���2'n��y'g�t�A������tQ�p�"?�᎑H��{R'�kF�:Y������eW="����f�v�i�Oz��QK���T9�.���^]��?��;��e�%iX�bE�A����48R�S��C�@�
}t����������	�<n(�˟`p)�7��$u�cF�[)*�D�o��H��c�Wtp,
����S�[">���f�y��7�/T��Ɖ�D_�Ke���<
}�Zɨg�#X��p����$�e?,�����d�q��愅����ՔuN��ѓ�����S�~:��=B:8���w�CΟl��5��`��`�@��Te�wC���X��a]��	w�:��V��8ؙ�(x�D��Ec��B^�+��:_x��9aȋ�	��I�6�:"wA�)m}:c%��	͹3n[�V~�Z.A)�������^�ﵢ�t�*2B�&�͔w\��J��wU|�*�P%-(֭N�֥o�7���R��(�rx��Y���2�G�3��_�C�
� ��ǲR�uƦ�C��Ξ������5�a� 9��_��q���K�C����Z�u����d(�u ཹ8���C9��W�_��gO�3E)2���U�o'\9����[���[9`/���|��y��2�'.X����V�W��i�7sH�t�3����uJɴ�В��0Y���
�L�aQryHE@�V�0Lm�ш�;�E��'q�8��h���ݜ0��~S�SQ��l(�i���9�$�RפŽ���m�!��/1 ��UT7��\4���r��W�4�!�*�ܕ
٨
��H����L<%E�.H��	r���Ld����s!b�l�UD؟&��N�Dź�ن�r���yH)�@0�'^�b����_,��U���U;� �>�u��͘�g;�ɮT@����Ņ�����X�F�5Dy粜�����|��[l0��=n/�᷵m<����6��/���r��80�͙`�؝5r,��j�=@��GNc���f^]�pV���)p�ʋ��B�l	��إ�-��h`[% *YC��h	�ذn6Jw�0ui�ꆼ�+ccը?U�����ò�j��y�-�s�z,��ָ'��7������D��x�ΡN8�6�#�x�ƣq۾��ޒ��M��<U/�s䐺��eSY���T1��s'E<@+�G��f�JD�A=���?�Y�\ӑ�F0F���d��g�p�2,gx���3h
Չs�$-�|���[]����`���h��J��kZ��W�d4]kՠ�i�n�l���-NŦ���H�2����}#�s�[G�8�C���&������>��Svg�P�0dBy�,�?���K�0� �([@c'׊�Uj�/��@� YZ���׽�y��Ĩ�Z��S�-(ghu]�0WO3�&�a�yTX�HW`=i��S�EK�=��n�/�YU|��2H���q��X�O/Bc)�
8;v��'_XY�#���n�'5�H��.��LM����6@�[��C�Pz1�V�^�䘩���H�b}S��9�Gl
1c`=���.;��/�����I�Zx�L0�.��M�6�� Y�s]��,C�%oeM���>b3�� �������po�=-{�oAK���e3��0,���篹��T�;�A�Wi���^	%�[�������a� TlHZZx��`S�'w���_�7'@�������&�z��yGX���e$���1v��.��Mx���0��D�7g�\�j���O���,�H8�8��3ڻ�o���3�k���JT�Uf�L�Y/�F�J�%��� � �{��Q7�w���ђ���	� ���������/usy磻��cDH����/��B��xl��O ��Wxr���D�|���Yi���2ؙU���o��dvJ�u���H�I�g)���CC�#���/� ���z���'�E�D����׀���lݱ�$�C^�q�����������W���0��h�7�㮯�jm���<A�G˲a����H
dZ[�߮2ė�Ч�K��ё�&c�����B��F��s� �\��R�`� QQ��Gh�/�����Ζ��Mn +�e3]C��p���(B� �[=���2�Xy�^y\C����ǉM��g��Ȋޔ���0��f9RN'�n$݆��j-�fƂ呧�"|�Ds�H����UK)�mV��j�W~����́s�i�t�X����j���"���Ƴ6���*� ;�%�0� �Gtlk��q*S�kg���V0!Iocdl�{�	�A���{����!������#-���$n
��}䊇*d7�C�EE��_@�\cly�f�+#ȣGB�J�Fv���`�+�{_�e�%>�s������J�Hm�^��x^[G�r�Y�ql�/F��7��գ�@P��22V���б�F�n��i!�*$0,uE����:>fA~9^ݼf#��r�HW�IC�(�K���˳5̬y+f	�3���S{�JK�k屇#T�3{�)EXG�8������c!�-H?ٵw�^�!s2�����?�����X5L~:��N�ī��C�P�|���>C�kՅ�_�	���OԐJ�1�+M��҂^S�uϖ���u�'Cֈ}�Ķ ��'C��O5"�w���� �_! �Z6Kט6��F�
ϴ�c6Y��8 L&�Cx1|4&$,pb����^�ל+��y�}��������g�ǜe$�_���ދ�E�`I��(��#~�lTu~��Lf�o 8��\���D�d�%%D�g:��!�Ed�4���sZs�X��@����A�c�-�����N·:��:� �5k�Ӏa�w��Yp�8*�0��k��4��s�_3Z����BE�B�^�;X�9����b�!@�d��ܺ��s+���l%�A"S�����V��,�{F_L D�1����h�Z��;�]����ۨN-���@���Tt k�7m4�����>�����6��ϒ�h��p���-O/t?�h3���Ww���z�Zy��t�� ��6b璨>�a��X��'m��p��������<7�cJ�QwC�N-��'y�TK���n�w�~��Ai�D	5˘J��-h�l�"s�C�doؼ�J�.��s/�'�ߺ��K�\�*�N��bӤ�&sU"�Jݹ�#L��H��-�zC��n�yW1�@��)	Dܐ����n�\R�_x?�y� K�9J>�hs׸Z�}�w����1X=�����8�]�� �;]c9K��A�O���|��K�=�O�H����k�-��{���}�G�M���d����G|N�y�g�&�Έ��E3��Y������>�_<�����4E��'+��8J��ȶ1Y��f�!�o������w�EnX^�A؆w���c��%�n�Q���Hw�Г�B[��yKZ������-��K�4�p����q�G� ���U���ʈn����M���}	���l+@�h�������G�H;U��:�8�ߙ1�}��nD��i)�9�E�uT-��7����$5�-͈*�H���7]��Qy���/h@�l׎�IN�e�2���|zc��0���ӊ���O?��
�N�e
�3�j�(K�	5�Q؀O�EP�y7M�Nݣ�ڂt���Y���D��]6k��b,�/��Z��������$�94u%������o3_�D���
��I7j�ё�c(���޽�*C[���4��ˉ6@lXQR9�5�zl����k�ْ�I rZ��F�yJ~M�{��l� H���4�1��9��������ӓ��+0`z.u���[L. �j�ǂ4t�9Z�մ�M_d�����\|�&1�z�w$�ȹl̓eP99R��^JA���w +���_�Z���f߈���S�ܧV%���~�.��59� ԱL���j;���^yRVä]���v�4q�r[f��s�(x��d#;<>x��眡Ц�\�x���?�Z=��a`��(�W@H��%Z��W��S�L��H��~�e���8X����8Q+�H����B�������?��&��.R���$V[/Z�Ns�����#9;��i�DȠ��{�zdf���t�{�g��u�U�XlУ��j5{f�䅍�r>-t����a�B�w=�Lj�C����j�e��H����BzS[�:J!_N���v�Y����g�e����*����k �/��� R&�ʨq�����+�����ܲzY� >�/�I�I�)N���B����]>(}�-۴�ʘ�I߉ڼ�	�.~��y
����xCW��9�ԡ�W�nx�NhgbDꗺ�\�G�����/ĥ0�fiyUBm0�e�6���3^���/<�8l����ʰu�X�"Rs�G-�R��*G��(�~p\�r�@�\���/�R����7�U&G~SO����+�2]K���h�O��gz<^<�δ:�i^7�7���'8��׽��u�5<�cY6RZ�uJ��,�/}n��Ļ�4��yfƷ9�<4a̟�����X2��Ҋ���sOz_T�?�n�D[f�iREC�Z�7�����dx���ݛW��Y�7C%��x/XL�������s���Rj_��|2DNw�'A,�Ű2�P���zF����	�@@o��! �R'q�l�ٌِ�����#��3���Tq�~\� |��Lj܀�%��s�MRL�鯛WL��b�����E�@R���S���G��k���r��.��5�rU��y�Oq1�=F3WN&����j���@dTN��N9�3[߰I,������Ɏ�Ե=z��A�$n�@<Ĕ*����$t䢱T�%�2�n0�Е�Z
D��QW53A�xId�I:�8�p�q<s�G�F�r�l��;�?��|�F�W�ZU���g�4_�|u��������^r��hCJ���i�	RckHc���]��N�v��o��-��7����!�\t���9؟�ʥ.��)80�Ø������YsA��������t�ƨ��8��Wm���W�|}�$�� A�I7�Tu�cW�K#�#;�!msz+P�R!+�s�"�+���+��}�nv����=��)��bb�5������_Y���#���ti��l<�:��G��23(�[����;=���HA�"�3�o�w�.��������uF�����L������I>�jsnZ:z�]g��X��l���:�Z�#�xk��'WO�0�$�3,�$lh1XO�����@+��wz�9�^�O7��;@��eX�S'�W���G�O�X�:�D�LO��
��&*N�Q�h�ʶ�]��o��-ަ���@|(�B/�ZC�k֒5�;M)x���S������1��*�bt2��4VY�HcΎ��}HO2��0��.1�վ��f�5��*�%�y�G����^���M���'a���8�� ��'�ϦIо��]��U�=�?9�߼�C�ɺU���
�z�@�{r�����~j��k��> �J理�C�-��,r�#��+(H��Ѝ#ͧ3K3m�:)6E���0�08\g��׀���X�D���E���p�Pu��V[�L��gv�+7�ud��A*H�"��c5��2������Y��&�U����-㿉پi�^L�+��Vs�+��]����zY9�s`6��Ƹ�W}�8�Gx{��]Z�#5��8"��ځ!&��b@�B��o}��Se&�=�!&�"�d=�,Eκ��j̳�n�dԞp��8%�8������ى�tlXU1����ޕ��K/J��t��T*���*ڥ�D�6�$z�Lg?�;cl@�� �k��u���=5�3���V��2-@�G�0���\FQ'}š�Qa�B��6�=�̝��2]���?`[p�N�{�G�,��>d��I���V����aLc
��^z�ï�tT���*�hX$e̃�� 0B��7�`�f�5+D5z�b�:Ҡ���ڣ�Z�j����ś�,#�h#�K�C"�����ӈ�,��u�t�� 冤�.7�脺��Yh���|S��,��8KW-�ӈĠ/��H&U֫���a��m��0��A��������ZRM����ҦL���Xʎ���7��Y)� 8i�#P�!�Ɯ�e*	���_�*���p	7t20��b$u�KO5�x�g�@l^w�<�L�`�:��I������>���%�O�,pwb%ԧI��S |mp�Z�)�%�
�=.8?$�J�i[��Gڱ`^F�����A���Y��a�E���|��6�R�l�v��cӢ;�I�5vF`�s(d>�|�j���,��4ӝ��}/����	(t�(h�F�����ZԦ��D���������߆�]ًjeYJ��sH	.N�;uL�է�7-kà����BS��#��4�6b��ϡ4��Z�2!KE(ZrSy�D
��d y]S$�.�X��y~�-n҆L��QX��U������
�����'�'���k;�V��~t-B�	GnI�'�?ۤB&��|��\p�pN&uB�a(p� ��AM����֫h~u\��?�/�r��W�c�� �6�l�l�ⵊ���kH������I�sЎF�W�5��L�v�b��{�����{#�8����T��۬6-�s�!�r0�������0��5XN j����NJ�O���]�2od��iG�����m�i��
]xOS$�i���������_8�@$Fϔ֔��T;p��O10k�Э���{�P2�
��L�����s�-�� �i}I8_���V�@I�7H׋�?�b�z訿N�v1���VQ%� �gJ1��<�H�C�j�2��s���9��	�Gj�i�|�t��A�Ѵ������B}񟞭�E��ˡ�v��p�M0�k��p)�s�1��e�A�x ����6�5j�MղAJ����@�)=��?�1�*�6�Q�͗C©�h�v)����;<���>4�f��M���P����3�+}�y��ˑ�ć���ף�a�|i�	c2��H�
��\��/i��M@@����i�;|��㸁���$�H��؞�����2%���^Q�}���Jњ��ڥvOdY���Օg9�Q�#��9�4M�A�I���+�|���1!;v�l+�������TM��3h ��n�7�~y�����f���H ݅�`�
.I�H�/y'�&م�DY�vt:-��wT���*����2m���B�Q��n�sA��)�64���fYK}��c߹l�˨[T봼%�,~�Ż��l,)o�u�����(�����\�h��c����F_�0��l��4эEB�mB� G)�G�L�[~�NJ�9��L/��WF{SNLVP�K�ӊ��;�B:�.<���6Y�"�I{�+L8U!,�TM%%����r��e<d��kU�#�k��Ժ!�E���m�<��)��v����u����*�詢��P��Hr:��^{d�U�>G	����+�l������uZNYM�K�1,|3B��;+�P�6�Y�����F�O��)��pA2���(��VN'W�(\�����&���4�*Q��X��јQ2J�|+��
n'z$�9EM$��)�hz�� f�`�\��\�����3޺Y�	�+���=� �t1�R����k��}qLc� �X?Qs�Un��rP��:Ic�8����̐��c�H_|e֛�α#v�@�eA�(V����e�[�!9�"h�vg���d����/#w�T�W������`��Y)�N+����
G;��E���D�T�J!VW9v�I�߻�;��hVC��x9LQ��%.2w��2���4�z��:5?q��'�~<E�[=��ꥅ��s]Ew���a���T�����{��a����:�u�J��%FB�ˇ	�4��Q�����L�z~��#?�LS���=N�xO�ȣ�c? ���]O�w�H:N|s�^�M�f���l~[�Ey��XE,�N�$����|�.�N�q����4���@�������8H7<����iu�?�i�<����P䅜>�D~���R���x�(EB4�.Q�Er�Js��G����N��ݨN����S���_��������Bga�ޖB����NH�E�d�*��
Y�! �,��Z�b7 �m��� ���m�y�O��2m2�S�h�xo���F#�K`���W�F�y]\�%6.��x1�t�C#���u���`�:�-���	����$b)��^ ��l�q`I��Ah���k�:d���ɏeR�l�=�N�tO/IE?�x:ʅO�`�Y�CEkKH�ל��k5��c������Ӹ'uEL�k8_>5R�Zn͝�/�]zcS�-��GC����x`��s�@��Xv�a�"�@u�����F[�7f�ϱڒ[Bz�%���̓�JWׇ�T��M��!!]�n�\vB�i8Ν���q�J�+�G���{��}�2�X���^g���^���%�����"̨U���WŊ.�n�����%<�ڟ�nB��ܖX,C�N���C:��:�.g�2@B�H�4^���a���%�\����Ot �Ѕ0B��"�/};�Tt-���{~w<��C8���,Ț�6���]yG�Jw�w�$I���nI��2^�W�Ϭǲ$y��ox1����;N�d��;� ���Вs.��	}ʄ�\����!е��<ٙ;]�{���\��b#ԃ��u�s�2e7�K�lz�B��.��EG}�����0B��c�S.t�Gq�i��_��>����Ay}�؁����J�'鿀%"�j�>$�)/.�k�X�A,oʡ���GUt��6�ެÞ�-[�w,n��ġ���]���+~���⫋�ZV��\!��0����DE"�m��Oݺt�E58��O��Ŷ{�!^�z7���)���6�[�oRw��_�n?�:���r��3�B����< �Tm��ݞ�ةL-{&�T����M}AXP-��M�M�]��?zZ��@���e�����������!޸�8�|:���x/���z��l�0�M�i�,�ڲO�Y�G���Ã\�'SLj�059�m-��.
ǡU!��k��ٴ��p�z��5.�B	\HC���u�UF��fl�������8hͽ��vcr�pq�r}s1��s~3d&u��Z4��mr�ڢ"�TSm^8ę64��󋁁Pu���/�=J*�>�������N�٣��@����c�E2v�E�:��Y����4>�����Q^hӎ0ig;�h3%~\�`�y�<h��B�_V�����R���Ԗ�U�̐�6~��^�P��ܳ�� ���@�����0�F����@���R�B�Z�E�����]onQ����Y�*G��_�Z��H�Zj26�$'O���3Mo���qy�L~	�� �ي�o0�k �y���]��?��q�
�_%�U�q	�)(���Ӫ�Y&{��
x���N��G˨���~q)�:T�Zׇkj|�|�W�ā~�J�k|:gȿ��V �Sɫ����_^r/>XX��)���5�TI=�3�?�����N��L�&$��;����T8�T���e,H�o�W'�Xfw���jt<�OQ*sMG߿����З�Q=j@.�.%M� PrbA�����@,��IzG�?�����jtM�M�����+��-=�����b�Qm�"'�¸T�e+Gr��1=��0g� U�n0�i�/�a�s�"��vs�74toFz�uNp�B���Na��5�9�)����~���)���Blt��Ռ ��*������~�`�%.Ec�x�
��v؅p/6#��&�G��uǟxpd�m��O �ѧI�qv��|z���v�W.g$sz��!ſ�@Y"HӤ�77\�bo~��O{`㴾����=N�Ƒ�l&��;��O���U0H=�-����$�r�[_8|eO���u��7��W����kiɖ���x
}�#�'��^DuJԇt�v�e �k��^�X�'�Q�Y�b��vT���Q�9���E��\��&@��G��vj^I8�\>�_�ddF�/A}�����J��L�[�����c���V�n��O���J���A��"����Ȝ�����-�ፄjh���3%�9�"����D¸,��w�9�ͥ�5�`�em�v��b��69����N[&K�7M�������c�5P?0�e٘<�h2WN���4�ӃW>%`� �qmB���9�ĵ<�J�q��i�敉�kxc���$�v<�Pl%���bo+#�{7v��G��:��c��Ν��wH��]�𴪶��٪��4���xrS���+t��R�5��]�θ ����u��mNd���W-��d���]�f�B�$��������*��E�b�fU�/7"vC�ڴ��[ѹt�7vJ�T�m�8a�ŉ�����(ı#KJ(��Z�}(̞<�`��0�p���26]�=)���R��GM�X�<�� r��Mf̏'�.�'�U���:�3n�jP�(�F�c����y�6k����?"<#X�O�g��"���4 \��p��`R(������/'��t��V�c�	JWD���
��v ˿:z]�3!^���*�J���Kh�R�׼����8��4lٳ"��l@΃r�x�[.`�i��h^ˋ�p�q��)�E�:x�.�t�G%�ϻ�jm�HIi ��1+͙T�b��Gv�=�,`�2%�q���\SJ�>_���<��8rt�_���A�p��Xd��51�x_�ON�ir�b�Y�.q\��r��&�]�M�J�CǓdDsW-݆� fd��z�#c��-~�B��"M�L[^�ο�ͤ�2@���=>V�l
X{��n��-���d��|��4A�U	��Ϳ\���.�I|#�,�F��6����F����u�yS��n�!wR��	Ю2M|Gk9�2`>�FX��=�Q�x��h�6͆��,�hf��3dｑ�7B-�i1g%�U�~�O���&����hD�XH��>B��S�9?_��<�>�ۂT�aFz��R�1Sp��E���$�!�?Q��iux��3ֳ0<���7��o�5ު��,ɒ0�D�ɢ�T'�٘��8�F��]����P$��c�4��=���:�c�j���?K�vf$<U����o����)z� $�U�e&E��έ����ַ{ ��FE� F=��?d~�aM/;�,U'�L�"o�(u�U2/"���8q�Ȕ��Rg&��	g٫Ϯ�1��2�"DߌL��j�f=.�n�cuw��b$��� P�zs�^��7 ֞#c9�ǹ��U'�$'�����Ρ��Z�3}XZ2��_?t�s�o�� �7��X���#��9�����GJs�t�hŵ}zVz8�0�xG� ����Ʌ���t�s���ɟzܽ�݌��9��	� ��"�k�$��������VhcnIy�<��`��c�k[G�x��9�� ������d*W��u�e��0'ʣ?r���gԅ���r��-V�2�	�pJ����3��ր�#FCb'�o����Ciy��i�jp�M�����R��VV�;�=.��7o���;en����|=J�Jk���Yw-�쐖'f�]^��4��nN����qe:��
�^Yh_k��U�m�?�4L��I�3���4�w')�v�b& ���x+p?^p�!���E5�)�~��� ZV~pc�9�Oܑ�D����ૃ����>���I�
r0�آ�K���y9��O��"�s�t+��,�=8ݲ�(��opI�W�]ǒ�v!����p�M�@/-^�b֖�i��3r����
=�b�Q���h#_�� ����\���}��+tG?-dї��'SL����|�Z�WW&�c2T"��mJ*̖\я5�����|��E0��M⑀��o�P�5�/'�5ЋO''��S�j��;7�ɱ	1p�$$Лp4o.�����¡u����|���v)y�)��.�F߯<�y=��Q�=��ez˃���rJ�'2I���<w�����nS���%B%��#M���}$%��]r(8e�Qaq����1RI��wYIQ���,H��Jdb�r�$���xn���o���z��=����TK2� �A�My���y�7��Š��rP��>ۣ��n��P�=�h�t��n���5zĲY�Y�/�GYZ��J�����i:���L���$�Nɀ�%�W&'ݸ>˖:��mG���Di�uؚ��x5��}�X/�k~cp��#��s�0g�e�C��34�X����9"R�+N~�+�`m�c��īV<�u��9�2B�B��q���	�n���og^��	`w�O�Bq��!�Aj�9Ⱦ�ML�,B�B*���k�ɀ�+����T��HMӟ8�q$���#	��}��X>쵠%����u̫�]ڕ>��=0W�@ȘH�8�T��j ��A�(��(������i��e�Ѿ'�˄��Jp���V�X��\L�K�������ӣ��0��[g�}�Qi��J1�����4��R�f���aw���������6d��X��h���X�n�nya6���u4�3���_�$�M5e����K��9��~o�-�A�bD��q.#��ݿ�q�����F���|\1�؊@��>y^�\.���DK��Q�R�@����A:��`����.���讆���0Fe�S�����g�B#)����-r"�!�e���lJ�9,�F*��r��D�;0q<��5�%a(j$x2|�q�a��PO��ǭu��B��:oŕ��z����WA��������;�Y.��J����v�i,�7:�$���۽���2;���#�VO����Gi�����C�h��du�)$�	*tj˼R���>�:�Jv��e���,����</��/۠
�ǹo�R.��,�*2�!��jG���^e9��W����ɣQ6[E��R4�ҍ&���g�4��=o�H�ZٻO��W���3S[C���B=��r9���;��2,ڂ�L�{Y�1�f�p�5�r���Uv����aF����jƞ�|����I��T�+�'��@	;
.o�B�g���
�)"�[��/3,pgD"�3�Z���i�iG_0E51 m8����uՇ�(m���
TܱB<"	���/��kt��4U-L9�-kxMǰ���4�2x�rC��S�8y9���Q"RNY�w�F:\	�VY��u��L�[���Ƌ�қo��Jt�Jg\��:"�PU��� �A�L �[!5��f�t?��=;XY0Y�Ѓ2!B�(�qY��T� 
�?N�~�u���=@�D�6�1������O�u�6E�Ν�������#t�������:��+!��ۜR����qf�%�BE?�o�8E��A9�MP?Sگ��Aux��[o�?��{A�3�ƅm�k���Y�#��(�	U��āC�M��&Kk��jnNӇ!�4�0�zx�E����TC�j�C�#:��[}���F͍�<�`����%*��㲻/�*��>�ǠȞ!!�����¿�	�5U�~?�l�)���	� RǏI`2%2�����ZSIg�qňYUs��d]�ӱ3sɾ�1�Ʉ#�����v�'�>Za���$�ݰ�:w�L����
��!�c�`�Pduۆ���S�h�5�-u��z\�&�gq/�tN�����cU3Ֆ�]�<[<1�껿��A���K�XM�l�n�6���G}�ݣ���_4�aX���N�\�cn�EG��op��XM�5����I�	��G����Y�Љk�Q�����*E��*�kq5d�^(���^rʿ��t�d��[�z���?����<�|��("��1���l�v�AP���<�^�>>$,�(�I����Rg�<��0�E^����"��n~u��w4��dЯ'W���ts}_��`��2h�Y_��8 �%�
e	���y7ҢN�&�ڗ<������x�N�l5�����Bµ Ԓ?XR:�������L���#�'fF?�����*� ����Ƅ&ۈX~tG�v���*c���Qup"aǺ���'K2���N��-�8d�Q�R�����m��"�=�x<�UEM�z�!�A`]���7�Wͯ��+��qH��y8
����N�9$	f���NX�[��1�����-6�>~�Ld���l>�1 9�$JϤ�2+�S��7�����R���x|������G}O�5T5�G]���GPR��/��'���rXM�^�������rQ3�t�M��/1�C;��c�z�[�OI�/]�]����#�(E��E@^o@�U��`�]���|
�2�
r����3K�։D��?e��qs[�,l8���I'g!����Q��#�3�����b9�s](8�X�?��>�I�XH����D�d����� �*h�`"b"6@��IA:���Z�_��D�d�����#��X�CwUoRdᝧu+�@��9)���W�iyG��w��{�T�OQ�E�������w�i��s�� o��l�1�^E�59��S�7ٲ�O{p�^عD5�ɳ)�����q����^�#���gε�v�?���bk�NPTe�]�$�ٟ��l圞�$^X݀-��"6���N��`Ď2�����h��0���AEl�,^�P�BE-�,�/��� �D��@�R�Ja�<LM�QL�^�K�z�Au����j,́b�X��0q4i*�?���Vle9�y��ݹ�� �Xvj����$�l���E�j�o"*o3��~^D�2���%�z걣 ���C�rᨘ��MV9��C7Ok^(�<I����δ2��Q�D��׉qx��I�[��T�@����\{g�o=��h�����}�5�U{?dz�o@Z� �H�徫��3��J��:�g�|���>R�6��W��.��������]l����B��&��
܇JgRӚ�,��z���'�4	���9D��II�O#���c-/&��C�>��jv��YM��/HHF�i_7�hy�qIۺ<Eс$fo6</&Q�vO�tN�t�cJCA�"~�z4qkb��,�`Ƣ	-��eL��9�Y=�O���Z)'��ӣih�'4�a���A <�ˆ���d��_؃��]��=��՟�}��-��[��jF�r004��s"�����׸*CͶLA� ޹#6C�pj�]'kj-�+�0v��#=��y?2a^+
V�a��K��ʙ���&� 8��x�o^]�4�b��E�ր��,
�͌�p��ӳL�{<t0����yt����t�-Q���W�-i�5����eP<�T�Iid Ȑ�V~��>�������rIIl�%3�%�.����3!��R�n����u��u��oS��ʾ�BZ�^��'������u�U�����dLY���j{̴k��H�,�N���A�>��4��0���=C��|���4�>��>�1����j�����f��_���~K�$̼;`�`[}0�	U���$ ��y`�eP�g:�ŐQ$��k�
���EN�(��~#���y�>��&��]S��k=(0#�Pg5T�Mܐa�8�fj �=Q�;����=@�xi�Z������t=�},�woTM��z��L�֡5��ܮ�"��>���!�-t�f��o<bA�ף��f2L�g��9�f���E9/פ�@���|����5����q�R�gė�k��f� UU��1��OQ~V)4M�S��`+��5otԂñ���$^��lót��q�k!n�]�&�/��6L[��Ƈ���w6�u(�'d;�@���dG={�1E���s�;�*�J�)�%Y�k�2-]��Ö'����]S�.8j,�;�:�yI^qԴ]�*���x����wb2{^}AޯiV��h��r�\ﹽ�# �	U��R�8�A��"�6�tS|��I���3wQ?��d��d��Y�c��S�A}1��[� ����y(��;��j��(|�m���(gd�x��ࡲ!��ŵv���:����L��YD�KEܮ �C����O�� �]�#�L� 4�l�,��^��.���6�@DCMq����}�)��͎q�j1�0�'K{M�wlGQf}/u�z=*ć{�R�)!j]�q�&�׸�N5�ӥ�_�\R��	e�y,��[sTZA^�+��8�����ǉ�6rr&�����SQ�{�Ql/Ë��#�(#Kv��q����q�R_gʶ����9�H-��r�&:.���)8�q� g�NRM0�C��P13�3�������z��0G6�u�0H�#Н�!���̗Qb^J��:Y�؍���U�÷hPs�E��g\	=���J����޷ù��vϽd5���tq���}¿Rr!%��Аz���]T�kI��˛U�p%�����_U~�,���z���ٶd�#��r*K����Ci^¯u����B�`�+k�M�+�[Ɖ��{���f�H)1�����F�W����Vq�q�23��m������i��KR&%�bv8�`��z��Մ�vW�O��;fN�j�6R��lp͍_rSF����(�ö���}�t�=`�m�=s��ˠ�f��0��Ö�o�sZ��E���0��Fd�䏲�`X�{&�����?sÓ@2���#p�p��x@!ϖ�z���Q�#�;{M��o{�����<:g��&+ <b2x`���дi�  Z$dLf�����gqS��,'F�(�{���Ҧ��k6%����/=�~SI�D��_�w��:�"!q�[q��tT�=3Ūf��H�s[Y[4 +"K|���f,�/���B~�U㯬�ц��Dk���|�o�/b�K9|s�Z�,��Ɨ���"��W��Av�����ߡ@i�$�n�k�V�^���@���!�Ç���e�:�"+صu���?�<a ���e��ߐjՙ������2�rj	���*�N�VWmġZ	UXa�5|�A��8^��Z���q"]��;>V4�s�#�i��;�����~0����o`�ТqlKY�??6ޔ|�	�������~�*iB�\�?q����ֹ=����1�-�~���v�1�<u���uN���k�:����d�ۚ��h�$4u�AƩs�dG=M��cMT�i#��xO���r�Nn�|��8��,��b�Lŕ�Մ)��q�@��2�*v�!� q�U�r���Z��<V���;������H<��ŻSD��m�S���%��ἄ+%����G2���։F1ɐ��:���= ���/rMTǿ_�?#G	�`��m�8�r�E�Il��8��g��d.��������A�1�V^��K-)H����S��и��!=�Q��W��6�f�P��h��(kc�2��A�X���͏�� /f�$hg	mIK�����(DŌx=��ܾ%k��`X�"a�z/1�[�\Kj�����He��G���]}|?�Fb~�����M�+�-
�!,���_G^�b����IK:mn@��57���-��2����m����quu��m����Q�=pv#F�q��Td���X&�l���K~u4x�iW�%�����	���6%���[渴C-��6�g|����M�D�oj/� ���(�:��gm)��.�p����@Pƙ&�Jꃆ	t��)M?1������Z�j�f�2W҉��������r�|��̓ğs��oh����j��ĳ�g��RVh�H�A!�s%*�ԭ�cY6�k��3��-Q����.�'OJm��Q4�!}'�����ߘ��[v���15~�J�`����Cw��Q>����?Cz˥�n_h����M�M$p���:l+kv�wm����&g�ܟ����䞘i򦦜ڰ��:_�kaL�	���{j�8N C,��?���e/�zD�����
>�$O���g�A%/�`�v.歆��w��Zz���Q��q�Ԃ����?�B� �!\Y`��_��h�z���h �ł�!j:�l���_e�A��_w�6�@���㛽����}��Є��M!U�Q�ow�#��5{խ��1�?[/W��TL3 �(�Ռ��#'~�E�i銚��	-rE?@��?��ȣc��%�Pd�Ĺ�y�qcp�z8�ȥ�$�:7H��ᕅ8�g/�Oe���
��$;q��<��d�����S�I֐���e1-X<*��^�-��o�1����D�Ϫ#)q������"�;��N#]b�|ɱ���vC�eا���i�"���)L-T���*˃Ї�)���6�$>ߜ��6�e���\齋��ԙ���P����s����<�䧗�j���A�|B�Zj5�<���uUi	��҃x9O����pV%6���%o� �#�把��Z��r��?D���n�=�K1Ќ>�Dz�W��� [�UL�F%|��畒��� "�׷��X�
�j���N�,ƛ5ej�m�5�y8R5��I����6���c��_���R4L M� Vr<#�-�(�{EV�Gݿ7w��E��2U�^�܎69����C�?L� d:4v�?�c.��sL̀���tt��jn�j~�OH�����6]��:Ô>t~B����Sz	�Dg�&�߷:3��X�,H���_k��F�n��/���ڨT$e
pg�`8H�:�wJu��	�v��?&���~�;
�෿/�Sդ��Ci�SU�"�'}X��A����K_ͮ�� �`��	��+�V�;e|���
�*>/��N�~I\��+��ej����o�#h��C���G	#>�v r	=q.�z\��K&.̔o�'� �^Y�5�x�OKtޥ
c��O�#�v(�B^v�UX��ƿH�}dъ����9�y��ҎɃ<��oG��˚�ȼ���(�\w,~O޴<�;�6�l4�t�/���!��b�)22	P�?4��"�4*Y�5����ݘ�ް��İ��Aa�<ޝ'A0Rg�����%p
�ǜ�G�p�s�w�*(�H����P�y*���'�-S�}������<�Q�yj$5���9CڔA@h`�j�"�D��O\�-�JL$�R=�Z�bi�&%F���q�̕z�)jC��R]��aLZ-���oآ<<�c�=�iS~��H����X��lb�ᮘ��u���:��f��Ó���m}��Uu���h����r�{�W��Ikg�^�{Gc$����C�K�5%Gy?rgk�a	Ү�����	&����� e,�(��*
N���TktLK;i��2
.�P�A�=b]�����2�c5��R��7���h�wǋ�&˹X�J��!T6a��5#~Ü.$!n^\L3V�G�� �Gt�/ƝwM��ʁ��:��j��ݍ�ߝ-G�זs��.���S�JN M����[0��:���<w�(&?،+�9�XGQ���n��-�F@@D���\C�U�%1�,����Y�� ��O�&����ן/��X34S��MR��,�nA����m�9{� ����� �⨝����؆9Lu�)���r�*��>i|�9<�'��J�V���I��ML�SQ���g���`/U޴r?Z�l���ɳ��t ?�M��:j�dr
������|�󡐂�0钝h=f��ƭ���)�b�g��
�*�?}�t^��xy�| �.��$�G�u�~�Wo=�J:�xtP��ስ=�i<�)g�c�����I�Z4U������-nX ���Iӌ������n���U�m��!�w����=���r.{��q�U�>d�x7���en34�4|�J�c��j!��ht�Ԋ�!�(].��*S�5e�wL'�Ȯ�K/OM����'��`��TYNRo�8;�����qK���&}�����d�ӥ"a��v����[i�UN�Q�'��0�B�ҞϞ�'��2D�P#�nNX���S+3�JJE
�[��=J(�G\��8]�@J԰��X��!�����/�u��������ӷ%�͎_͊4}�j�6`G�X�y�p20,{��S��	��Q����%I���H?t�Q���\���!�z�����ܴ|�'6�B��L��-�*�\��p�9�;S�ä́�p�#Q���z7�Cnx6�����vBپ�=UCɒ�'�`�~�\a�Z�2Ev�!0�N�
?�L�?2l�/b��D����k��fr�u6��s��	�!)��G���;�_t��2�pcU9��^߸V#�;j���C��7��_c۩������𐓊�|ԥf�^P1zy��p���	Ѐ������5��WL'�2�&�9���nٽ�fF��v��=S+;�k���oP�`��?B�d���[R�-���>h�e��d�،�Lr(Qp��J���� ��T�	 �W(ʫG��{��� ��ʐ��a^"	��ݛ��ЎZ��BF��&~��L;���%�G�Ă��W݊l%�nq
�Yt��8NP���qmE�{r\󍀮���ը$�Xae<{ax���Ы�Y���`��IF�����pQ� "i����X��%̯��Y�ޢ�]k]K�4��@>J���t��X1[Ρ��=9��CIogB�<���&Z��m���>���1D�6u!��	��}�d��T(��
��1�O�P�й��sD�ԏW�d���~�K�C�%�*1(�7|��B����q�n���5Q^����pWy�G)�ʿ�e`.��d��!�y+��*~���$C�C��Xg/"�����Cn�?�MӬ��R��m�����}�TO H�l�i-� ��l�jh�DLO���!_�)(k���J�7X詃���v���m����aҺSn_�˯s�~9��Y�:gT����47��j�Y?b|ۧϓ��)�杌�tZadQ���Ĵ��)	��l͍>&���,%'R�q�m�_
{b�:	�F�6��X�:�W�����ERdY�Wǲ!�����ɰO?�<F���4�Ĳ�����;&�ӆ�eصn���B����0nA���|ꉐ�k�Ն��K��b\^���6�Q��u]��9͚��kҾ3�]�o�E�M�Q�K��~�Gw�\C������Y�ZP]-siり,*_ݬW4YS���$��LӒwI6�IPJn����Q��(��W�~@��%��'�FAҥ�=�ЧG�<�]dN��,�Fd5gX��3�S#�O�F\U�	�<˶E �L�S�x�k ��/��q	b��}����q��ϙY�8�+�K���S��� �����H;�`+�WF�n[���*�
1j��
��'qaN�f=� �����~��(-��B��"�����)��Y�"�q�����;��YCL��L��L´u����i�~-Fu�m܊G'
�j�GӬ:}�)L !�M[6�G�R+�F #qq�s���D]�Y��!�w�����|@��M���b�4bA��ϱ���>���,�0�a���	�c�_���;9��ȹy@iXq�bd��
;dҋMFAR���X�|D�tt<;�0y�Y�D�+tW7%�x߰a���dHop�����A��$�v�!o:�eM�Ꟗ�(�@��N�(.n�n��������9	�`��@_��y��`y�(�W�OiC��+�e��u)(������!�:=̹�\��3����yM�����ǎ����qE9�F7�E����R�Q�<-)��b�n⼉p^�x����X �|�{~]8�?iJy���l��j#��-�q�٧(!,=��Ž�hu�)��}C2����A��阕g�I�)BX}l:�ru�';�'���t�nd�����A%Qj��,j"UU��pL3��{�@Z�F�#��$_�U�{�a|+K��hhH�NЋ`������0����.@�X)��xD�����_���4�Xi!��(��ϕ�$ �J�G"��"G^��[�dl8���,�_A�/�a��v*��S�[��
���2`�.i^�eq`�v(Ur�c�<q��A�Sj���)2A(x;*`���3��nt��d���v�������wvP�J�j�U���;z�����`��&{PŘU[~E5�6���.-�˼���QMP��M�^������б�����^�P�X���u����KB�AR;�������Պ����j��6Eb�MJHte��녤��	;�A��7��(��= �U����ўW-�Q�QB�F�N���>A"�?�������f	p��τh/��X�gin�p�m��j��=R=���^��L�v�mΕ�UNj|�\�aI������Y��]��?dVu��2�E�R0�<O���D1��j��_��䂎�w�\��9�re�e�=W�^�rg-����c�Ʊ��,�\���8����<��iW|�ƹ��_%�+�SwD��n��[�K��SQ&0r�8�}�t�#���`���Ks:\��ӓL*��w��[�����#�G�o��z�ʱ��������rl�!������c��e\>T�^�������YФd�=������i�����S�2!@]�z�аV;�3�Uj��n�Ǘ\q����A���F�?��TL�bݐ"š����Ē��h �hF!��I]���� m�&ɖ~�����j��FϪZ5�T���|ᗋ(N��I�>�YSy���[N��Јt3eR�fN|s���4�� y���T�ք����� 3��{����+W�Q�����U��Kkq���	\쎣�,a��C�h�U8�a�Z1v E��'���X����~��hUD�*�Ӥ�\�&h���<��ned�4��f�V��/7Xt���{�f��o:�d���Y
�r��{Uֆ��H�|#�o�0q.����B�.��J
`Dv��E���%Z������ұf�2��io ��g���Ʋ*�Qk��36یZ��͈��CY�"�R�������������ڭ������x��� h�R�~�`ItKx5��X#���y���_ ��7a�J#��l�(9L�Ԓ˼�Mx~`Dw0p������p\�kMx6X���~�U�U�/pw���iX
n/�»�cȫ�B��g��\�id��@�#�TD�3�Vze����%���,���������_<iθ�=��������SO�d#x�VB}ԛ�ۦ����,�.�����y9���Lc�^d/�]\>��w�cJ-��6ȡ�٠H�C�����p3`(��U���͌X�o:QVY����~�+8TR@�x��ɑܜ�F�׷�����v�u�#�5�@��]�<���B�g���6���C��)��H���uO����i�����g�H�Vڗ��Y�;E�8�`� ݿZl$���O�������'2��W���OK$|�t�R��ʃ�=��	N�T�~�j��*��݋Q<�Е;!��S�U/W�َ�3�����PtfQ���$?��L7暏��/��Z������V��P'IHC��&"���y2��<�m�`�[ƙ�z��LJ�ÄR<��-�©ϓ�!&NXSӿ؀��Ǧ�"?�Hk�#Qr �i��>�b`�����LqM6j⢾rۈ"Ȱ#�M|Oأ��޼?���G.�F����TD0^�_�۟"��oCYa�yrOf�A+!�#�c��:^*��]fY��:�{8�����:�ڝӚ���*/�d\OC��t�hi-D�W1G��qђ5���h�S�IE�����P�+� ��6/��u ��U}����T���+��BN;\K���Oڂ��՜F-�����u�u���`�����V�ėKؓ�0���2����Yj��Q=7篗p�\�ʗ+��"ĕ�¯g�]��߉�[+��4���5�E�o5���)�+�P�(ޡ��Ɂ�A��h�C*=��i��6�b���፼R$�9vI�J���$�!^6>��ɥ�}(�y!��fXi�9��Y��m}_���X���[+`��.OZ��t��X�ia
���tyF�>,��N����r
�g{�)�u������/E~�V�0L\f4�R%�fhY2b�W��hhk� ׅ�~	A�MX���
����9�X<��n��q�(��,�&��>e��E�^M�ѡ��0;�o�n�΁�Tj��9��0m�m�:���'�F���!߃26�vs�P�.(Ò�\^C�h��]m��h�l9�Sk��*V��T{���}Qi���2��i3i�cON�Ͽ�ej��C�N*��Y��Y�Y�3ЁF�8��0��Iިp�v��y&~��'�u�#qv�����S~8�ߞ�_��"Yo5���[��� ���xſ\��ڼ���MD���O{����ǔ�%��)w�K��k@��+_�#�q�ݻ6{6�#���i\�v�@�+2.*+���{^�	_L��0LNab�:�j�ڛ�[�F\%?1'$����*�C`#${������=�
�m���t�ߌ��np�ݕJ��~�Q�#;�X���7�#�*y(�܌Pv�ӣ3�j �hӄ�1�)k�q�Y�>�Pۭ���z&���|j����b���P��v;��[����GnYl2����6D���m�ڶ����ĺ�Yg.�8	Oaq�����>E�A�$Bw;�e��Y�;�=sɝݕ�V~ë�=�,
f�
ĕ�s�kYh"���3�F�IGMI<N{������
]�|���]D4�,%�wS"H�捌k���=NH����͓2���c�k4|��X��S�6C������8䁱��ת�ݦ�d���!ĭJB&$J�/�A�L��E�gTI^��$�*�)�	��3P5^(^jl����`|q�пы��0CZ�)�C��ŨV�^E��_b�&��_�u����]m�0M<!*�7��A1b���ܑ� L�b��[��� ��]P�Çަ;o��p*=�>4��7-�m&W1s:��̡���YV��A�n�i�����&�� ,���,�y��&��D)������b+��.{Btޡ�sk"�h�~��`�7P��3^6�L[����Lj�Ew��k��B��R�0�v剹�4��-���yJ�4�_l�@������=����޴{sKb���G�>�U)��4��	d\�k���~��2X��hl=�Q�d��W�ebh��/��q,)��K2lŶ� \B��D,�5Z"E��b,��'���R��@�R�6����?�)㨁���_��;S��	��~�cPiH9VCP�z����h/,�w9��"�yq+�8<�.	�Vѿ�s�����8O-2�8�3��;����9�*,�H����-�o�W6���eM[�ϩ��%\M�o�<����#XԘ;P�V`�q�  `&(�M�%FU�⛦��Xډ�&�ߏ�G����I���I����_�[]�c�Eȇ���&m�r���b*��;T��2F�v�C���%j`�:HR|p5�aP�T��Y�Jt�4�d�������,��<]~���DEߏ�xU>}��(�@:�aJ�咩R"�z�܀�T�ʏ= i�
�tԵ�9�3�����+�盂o�;�Kc1�F�N5c� �ȸ�j��_+�D#�[0%H3
�����9Ld^X���ƲU$�YDMbn�ڝ�
�<�~������I��ɗ��� -|=�e
���"*���y��G�%3_I1�h�(Wd&�#]��%�ʕ���p�h��A���m͙�gsQI���|XP�y���3���Y�&�cd�	.����or�n���X+ܮE7�-�0#B��Y��eu��g�Ҵ��8�������L��	ōo8G���&y�*W����By��U���t`bR��l8��4|�2�u��� e�Z)5�Z�˗�\q*��~
�/��f�:�2|��+t�4�@�T�N�� F�`=�E8�k�N׈0|��6� ��!N��9 �:�.�a3���i�tlnJ*�.����|�`�P�n%�\m�_1��a](�k4�
�Y�a��f��0MSj<�K��z$e��K��
͎N��5x��n���� R�ə��ͭBA/BV�ر�:V�׏鼂�xΊ��� ������[;�w��"�6��%S ,�;W��Q�!>S*��uw<��ij�奸A�Si��Ws���Q식3y��U�lL���'oʓ=�S�o5P�=���F�aPQ-��~ߒ�Ei�ӣ�w�AnS:x=�򋬈�!>��"N�R��ިA58q�	zu��ta�SL���'ᬶd��$a�~���+�$�
�Uk>/���l�g~.un��?�; 8��N.�X_o~�Fg��Ԣ�:�N�P��<��z�۩�裗�n�"Ɉ92�4>U�����8����:B�J/�c{i���/�YC��Lx�Ȏ}` xɢA�(C�`#�n�UP�D��*z�ݢ%��V�×����C+��g/�$60@w�~7�r'�,A�C���|ۧ�м�����r7e��Tw0q�7�%S�.�_~�F|3�#�80��0��I0�eHx���R������Z�̣�A�r�~ }h�D��Z	Kd}�Z�(�,�K�m�ߦ|��l|ag]P�g�6w-�R�Z�!�x\5U��M����sߑ~a��"+�Ç�L�|	�R��Ao�R�]JDT)_9���S����з�t�x)�n��o��n:��,�r�*��;�/�'��T\n~ø�e���j�����n�=\��ˑ5�[^�q�O�'Ë�*B�����$z����|'2��;&��="������l�,�6��So�c.&�z�LgX��ݡGj�~��6��im�j<�x��A��ID�j�w���2[�9�>+�B�`r<���+X���ަ�vpG���C욊����3��
�B\uǵK�b!� BO�z����EZ��Ntg��5����w��f{�zy�߃<� �C�@xm�>BqHl7Š���d��`��Y�2���߳�m����Fǐ���I��_nۋ/+�X)�cH�uh�ї6��BTK3����(c�:���M�*!]M�&`�k?�[_T�>J]n1�+y���斊bY�Ak�� ��m×8
��4��A�^��������CW"(��!=�dx��z�A-)�<\<rW_���1���j�Vm:8��z�{���ם@@PUHc٥+���n��Ǒ6ҘRu�*j��Th>Z^���@;�cf�+Cj��`P7i��iB��I.�F}-4k���2=./?f��BW�o�%IH��덂f�t����dg i �����S����ts{�q�E3yN�YC=O��Q]��s�$�K��0��I2R�6:�֫��@��6�L�S�P{|��k��ê���A��*8���cn�@�Qr
[@��#L�R㶰y}cD�l3>r�9"�5����j1�$,ɯBs5�V��� �=m�f2:.� ��6l�l�>11)W����Ƙwzr�����*c;/�y�	��dp>�@�F4�l�3��^vCW�!�m�%�9���7�[�5�y��6VݰاeIr�'���EbD��*:d-��-��T\�zc�� �7��aH9�\�i�w��gs���lW0�IH}�����7X������c�T��ƹ��H5�f�9;�d�<B@{K�ew%_ G��9��N,|��3"���v��H2) �I�4d8�����8	j��y�Y?U;ơ���ض�HJ�G����ޡTH�W{>��+�"���c�=|q	����{��=��@�@�V#�I�@jG>�젯Q��T����
r���!�3%�nֵ�NC���"�C�3�k�������>ܟ���������� ��ӭ h�=��#�K���<��9a���~	e�d�v��X� �N(k��5��\p(T=7R{�E��hz���|�g��*�D ��m�.��|/��]>:�RS����y<{�S6jqY �FG�E�J�j��Ň��lG�ޞ��(�b �s�>fn��꾗�����z���]�[jT�%ޖ!�I��u��g�V�[U��3�B��N�ʶQX��^{���_�>�L	�}�a<�L�rog�4�'����h�1��u혏@x���>ir[��4��kg�mp�`yt�d�|��e�$g2�Z�06�<�|���ƫ~ti�5E	�f
��A�M�4(@�"-c�$G*��#0�0��ӓ��&.djI�]V*ĵ{*���NJ�)��B�:����ċ[�	�w\)�_��p��D}��
/̆�����~�"�!�E
�HS��ߗ�f��"X����;.P����D�S����;K�FM�4�HUｲ�K�|��X| �L=��$#��wN)�����`�.����}�80�c`|_����n�q���Bq�aj۔�G.����ވ�1S)�` �6�VE6$f��k�NY�G��ز;Ks�~����X���t����ƽ��%�hq�\��?�*A�%�l����(�:3]�3vW���9]4����yO�Ih$F2]�_�=���[A��-�y��m����T|��d��ҶYϹ�ʘ�	��'Ѹ�T{�0z�x�f�S�����!m�[ �"D�DH[�GzR ��;��%�b[�#���6��m�w;I�n�g~C辁�2����A�Ƴ�����F`�-
�J'��tC��"�6�Qs�P����O�W��Kj'-{7$hmb��\VL�����Ԑ,L�l���g��.x�yy��+0Fx����U�a�������v�4�?U_��On���3������W��]�0z�!5��H���c�� �^ǟQs�:�6�h��X��'5��ߕo I�p�S�����ΐ���<H���j�n@T��~�����^SE�5������`���צ�����K�G�<yО
it�em����Lږ<sY�<�~��K�I�K��V���?��Q(I��X�Ɯ��A�9��J�1����e������[WJ��:.�	}�� ���\�K����Z9��p���G ��j�\���T~I������g�S���ֱ�HD=0�8p~�ʒ���R��D`�=�;Q��BXRK�D�����V�cZ�@ZJ��Fq�E��ί��j���Ԣ��|5�Q��b7i����_�Iʑ�H��<�tE��Γq�`,,2$	�U��;A�U��3��%ŝFRw��m$����d@�Ł�����c϶�C3����/�Xߍ�/�Q��=%�|}��>�m����R��&�J���Iu����0�OT��g�8	�������4�Xu�E��G��L��.P��O���/�F��l��׆JH�Y~H c�7�s�=sXc:��-���Nԑ���T�'�t���Ez�� |N�@�,O�"�׷3
�	�`�Iԗ&s���z�;z=}��+�a��Sw��i{�9?���A�
�6t�h)�u�3_*Z�{g�l���������i�U�%�U�ՠް����K$���ĳ&
t��˾na����{[�'0z�L����y3 L�.wF��R|�z��!S�q��� m�sϢ��bF2A�<��͑n�H?SQ����dǆg�k �6c'��8�¡��0~�ugGFb�/7>o���,m�)?�� ��5|��oX�6(�\5�e<j�Ö@�uxO]{���̠u�����ԟ�P)��ԥ�\������>����w�ʈdN�����P��������������V���k���laT(Q�ԙ���d�ˏ��>�]�b�b�S�i���K���!X��6*Dg�%����د$�9=��/~�{����vC���~N��7�:�����m��N�(~�@���`�d���g3�s�`#w��x�H��9�A(��7}B����L��(�fm)�l|��`S����p��q���Ýh���W�xC^�be�'��A�������
)bz�_��a��ܺ�2X=�eM����\��������\�kէ�҈Q���S��3�eu����Hc�C��9��/V^�_�����]�Ш�A�*��E �7�=�8,�ei����������i�و�.��`����˲���'P��]��T{�?�K����"�ħz�� T�E�ŶY5}�B��}#�Zhqv͋nK<%Xs{���gihf�IL��%��t(��:Gߕl�������芡j�{���<qss8#� ��Պ@�}dY���_t͠;�n�K��oH��>�u�$�7v��~����\�or;��z�"O��{�f�X?S��#�*��;/`�43�lȗF�d�����(^;+�3��d�pH �m�,z��id�#�4��p�RB"��:�	�]��NT�oo���q[H�nX	,E�i�~�+��
P @���3}G�	�f�A*n����떭<�H����D=ݺ�,3�VLQ��Hɤ�q�}��}��tm� a���Q&D�S�U\�Z�/go��|���ġԄ0�r�Z_��l�����_իP4{����'�eԭ�$�Zk�l^��ϼ��%
�#a���#�KȄ���>�m��\���zb+	Ӝ)v��Mߞ"��Ҭ�q`%���)��N`�F7ʻ�p>���3"�n��>B��M�Y�ā$�i�UI ��i�$�o]V�ߋ�ڼ�j5m,5���-�����Z���8&�!\k��C0�M݊��[�0bP������\�"�ܶ>1�49�ؕ
_"4���o۳��U4�?M;fp�o��؀yl�&!����wr����4��zjI4�c�J��:4���cR�\�����"�N�N�-;�Du9�f*M��� )ףC�C�U�ϴcމiƫ<�L	�m9���3�}*[}��g`A�:��]Ț�Ũ�G�;�������y|�>x�A%��P<��z|ߵavw%G9h������<���������_8ȗ��X���r))Ҭ�R���=X�sf�q��0f,t�e��KX�E�'-UO~<�yzQ��}z�f�1"d��ݰ~/,�ʫ�硫�>������G�,��ϭk��~5*rٺ��Պ��1~| �xc$�Ϊt8K��/ܤ�
8-Cv��\�t,m�͌��_�Es�qO�^yil� =�c�Ҏ.��,����>;ϛ��7��Ms�p�s!͟qk?E��A��1ig��6YZY���te7���&i��5�����i��I-�r1�đ{�&-o�f���6�s��QYHuG ~v_�����V������u�����$��O��x�pD��� �Ǩ�Y�`�_�@��Lvv�מn�z�j���� �CCdJ�i���]�1��}0��}"��|��<�E�l����B6�����v�����G�%�/�.^-��$�;im��%k;k��%"ׂ�HA�䟐/���[�k������	�e�X7f�^�a��B�ӗ���n+�+{5B��t��y��rh>)��ek�A~�M��v0ɥ6v@DV�Nl��2S�n��}�[P�P�~���&����+˓EwH^F����i�[�6`#%�~+��xK�[��Ҽg|�#��{�[�u�J\p� I�M�C%e���E�ۢc�!�a.L��.{4�;��W���|�$�=��Ѱ�8���@y����=�.�瘫��8��E\v�n��i���Dˉ������ONi[�Mdbɏ
5Y�G��6q�2�o�:ha�q��yN"����=�iֻ駾%�8^�oƸ�(&�]3o �.�xb���é�
�y}�=��l!�q\Wb��ӓi}2�%������fw5i�ڴI��k����4�#�
{�]���K��L� �� 	������zr���:���O�����NѯT�!���!{�R+��_�?ܭ���Vm�Ɲ���ڧ��&�fб1ѷ>���'�L9p�6�����Q���3h6�y�_���)<,2z���5�!H~�������
�� ��y]��;��@��q1��H%��r��b�[ƌz �s�Yaw���6h�u�MK���V�I���5��r#��@kV������ב�Q�#+��L
�m��5���N"ȧ[Z�r�@'����Y����������ۡ�t�ځ?�:��u�a�(��86jn*�e���bfBQtC0���i���d6u��k2dT��Ӳ&�U֮�62���U/MyQ�hv��-S/��d*+��FІ������,�N֤��:�YTTy1�(��p�7a1Q`�8�*�7:��'o	$�;�����3���9��
?S�Зny<��RD)�~�� R�Ȓ@���#tasΗ�CBk�x���5[���t�:9ꄁ��Ls�q��p�ZH�ó�j�c��K\��	�����\��FI�z���P��] ��[8ҿ)�G�H���h@�/Ad���M����i�ŏ��������F�SB�0���=�z�b��\|���M�M�i�*b��N�����b���k�6p^�=�d�y�^Ԛ�k��} 9�!�|v�4L� � ;�@��M��v����?c_�
�0ל�s�Uۅ�]�J�4
m$x�_����ʯ�3Ҧ(GnV��� �3�Ԋ��rq��&���i�_�	�ac�0�2pdΜX9J��'¾A�;a������u�^��Z��ّl-:�ڏ\���8���̗f��^���˪�Q˳d{���.�M�x3�v-�4`{���1�4�j2�� |�������ᵀ�L9�L�96J"Ϋ���ߕM�D[W۠T����E9�J�|Qr�_l,�/`�S�1똏�sNl+���T���:ƊQ���<1a�Z�(�p�d���@�w	b�:� ��ORǧ�� �hQh���js-��G���-.F>3�EJ��n�f�!,q� �����-Inaa�e!��9����:�%mіݵ	�� jiqϡ>l�	�|0@pmpX�O�T��{��e����J���o.����d��������}�V�EhִF��cH;������e�W��q���A������]w�jpù�!C�Z�~�VoA�|�`�{���ZY~�$�+�[M�Z]/M�&|�����F���\���u+��b })u��pv0�5����Z�w<+�_ ��s�^ �=&-�1!!�P�:�?�
���������X����)%���3�k��X�W~ر��`���;*��n�9{�}���5#�>�0�Q������P�wt������]>_]/	q��a�s��H�97�z��{�����Bc)Ӓ�'tf|Ҝ��7=�z�c��`����t&�w��#����6�9-G��.ߛN6����>ة]n���w4��1N~h��Bwkr/Fs_�e�C�J5�*��1iiu�zׂ��O�A=����̈Ԃ�Ѻ��xQ/I^��)~�c��t-�+�s�������,^��8�n��Ĭu��>ѡt�	<��C���>����
�N��}v�H<�nh�WQA��ߏ���%� ՞y���v�I�{��c�0�̩�?D��
���C)��*o5<�>��>@��K��S���t*�Z)�CÎt�5�;'��@`�O�4(RX
f�����ą��c�gl hl`*Wk���.O@�_�d���[�WL��z�5��r��S�F��φ���% �#�o����1���/���������S�D͕�gHvշ"���-9d�9�8`���������4L.�Mo��5�)j�0��e2W��' <ɬ�w�Wף(
]�'5!��/�����w�����lھ������D�^ɒ�� �j�$��~9�Be��.��5"`�C�-w�d��0�@��fA[��ޗxPYfX�7�C�<Қ�5���F�L&�H� ����Y>���߯8W�V��Ɠ����s]�B/5�Ve:lN�`��c����<M׏m�aK��(���������.��C(*����'L�|JRO0�\��LK�6t�^�d ��.���r��STי��'I @M�N��F��,F���MA, Þ�G��������в�Wnޥ�Y�:���>0ޡ�G{*�3~:���x�j]��,���*��En�qdզV���*�i-
-�[J2W����2t[�Pd���m
^�s�7!�qA��{��5$���-{�Z��X8J����%z�u��g�p��M����+�`�18H��x�2����3�!xL�;��B�m���*i�� F#L� s��vu�3�%��@L��j�K7'X���Q;.r ��lb��i��T�	��m�����J�w:��d�l��䮒���C�/k`����<qǦ&��V��w���u���~������Q{�<C�is���ʰ�	��V��I�JoA	n�Oa�/����c��d��_d��.g�R�5�u��Th���4 �X�l&��Kx�,�i��:!�XE�.������܊SiB	���x8+�a���<�&1�����2f�r������_�kk�|@�bnQݬk�mO6̯=�M�[��&���aP�Tiq����(��쟒dg8Л����í����ȍO�=Kܽ��Ea-�@B�;i�����~ԕ��7�۸�*���շF�9��fv�&W�p1Za��-nOOu����M�t#��]��Ae7ǓJ��
ed�bx�)�Ao�/�L��^􊇜'�E}Mt���U�_�l ?�%��UT�Q�h~�V �i휫��LG���>Z�q>�T�f�d&��»x��}�?v��_�Q�h���B�Im�ϝC��"��R�,�2��x[Ǉ��|ՠ���i�PH"M:�'�=��g(����>�*�R{ڐ�^VNcS>��2Ժ����w	��X{RwN�bp�a��hݜu,�>��e�P��y�������q��l`�JF'�N(��>���MB<q��S%?+�d�`z�t�m(eT�� ���s��ݜ5���ڬ쎉�ä�e����7�n�d�b�cI�̨�2e1�O�ևĺKɄѰ��ߜ��I���oq�es��Y	8!B��&ɶ�?�}��L�1�hZW7�67�t��\��1ٰ�K �'��ŧl�C�k�"�5���Z|S|P�^�+��L���Y�ȉ���&���)��$U�Ѓg������ m��[�̲?D]o�����%�J��z<�@؞�
4��&��]��(&��V��+���G`cҢ��b��$�|T��Vw��ڡ.��w����̏[K���n2��sGC`���W����}������7A��G��W��^,�Zح����{=_����D�f.߸���b�V�Z?�}3�v�oB!�t�q喋h�髍^!��˴�<2SO̖PX
�ۍ08J�>�"��-����J��������IY]r�!,�]�9#��l����k(KJ2�"�/�E�,�)uċk����!8X����yf����+����j�iɭp�CW��Pw�3xN)OW�dȀ�sm=�ӵ2�t@M���?��] �C���!�����/�|*Ӗ_e�ʽ;�ݽ�-6yi�K�Q �<t����ʑ~����'��,r>J�	[�����%���-Q��-J.W��~�
}�;<��;����2�"*��b��R8y��3�/�B�a3#�R�C�b�R�_�.Ы��K������z��b�>���ug�w���������V�H $t��(�
��D��ZxGc��GV���7	���8�1ڴ�4�	�w� �<6�����Ye2A	!H���-�K8f�)�t�ё ��`�x��hJ�]�#�t{k%���Ń\�>�{)��9����Ֆ��K��aU�]�j��,���q�,8VV�`K�,%��VP�{���n��g�VD<Z�×�=����h(c�>��|oI���l��S?D+}�>�������/�\"/F�PfC�}e5�y4I���s�x�6��(S��g���0Ø�����{��NK8m�UJ��Ҧ����څ�`�A@��8B�ʣ/�Ծ����n�L��w;i5C6vo�AGg����{���L��	�g��o�Ig���p�7�C��'J�|���*�_Ղk�P�-����˦�IB���ę�	�<��њ�4�l$T�$���q��:��o����B���%�r����qx
|n�qVZp'|�"�e�e@�q�6̟+��E@��ɚ*��R��.���P�Xp�o���%��)G���^4���)(\�i=�O(�~�Ϳѣ�d������x�1�!SÒ��f���R��-	�bOT<��=t�/�3]��޳H�fӥ!Mc#�f9���B�_�J���X���O
A���s���.YQm���m�6���-D���`�'��g1_�lʢL��h���f�@��}�fv�㛧c�[�����:]�W�k��E��cC	���pw䘮]X\X#�l�:_{����B/�r���ك����b_0R��&�A���z��u�0�c,�ק�Z�p���A�Jڙ����q��̎��Qn}^�գs�?���u�
��ق�nӧ33b�mk]�´�6l���!���+�$���[����y�qT҇I���l> K��R4Sv�R`FG��tP<z`k�0���o�)�����.X�#+"��pw1$�6!6J?���UBq�`���R��tI��p���1�z �!� D'��YjF���]�^�֢�EV-�=4�[H�+<���cG��A��!�G�)�Bq�����rZ��LT��
��P�TκG�!����a���Ty(y.�?([���<3���u8�ưn$�#������e������jM���+J.k 4+:�f�B����D��͕C�2
R�9.m�ny�b�� ���!�% %�PU�1�x�h��`ݞ��9�_�Gf��|�і��&��,��$5j�!�&��,ͩ U�)�<���î���89~`rP|��*�� ��ʦ,��(��b�#��n]9:�f��"�ɢb���A�L<�ZZq��!T'��-T)�D.P@���TYe�� 
;�bP�A�}�	�ymT3�B�I��z$�>�Cb]�ט�����|��<!���1�KY~[��K�5��H�n���VV�Q�R�
����3�p��K�SIW1�vf�@|f6��M��c��Aw���sXz1�k_6�w椔\f3D(|�ډ&�^������6b���A�B�����r�0����A����O�g�zGU��w�і�����0����C�.?����c�W>�Mqf̡�E�yw���;_��F��`�@����&Jf/�f�<�*���P~���)�2֗��6�R�2�D� ��BZ�����~|�>$(�&.�;O��YL�b ��w������*#�or;VtU����(O�s����0�H�ʐ�ƍD�1a�6ʈ
#f*�K��r�a�����vr�;ʑ���01O(ej������3���~W�����r9Y�>��bgx_���jY4Dm��H6W�̸S(����*�=H0:�@U�噪��Sڏsϗu���8ا�%wZ�� ���~�5���OתH�w��.yU#W�2[)�P*����X�Q�4ya
��frY��,LG�$�5u�r�p,���Fy[J�ee^m#5iuG��х�ǿY�uir�$�䐿?X<3�`���������}��fD5I��eJiO��Rk��E���T������q�DU�E
wh���H�AU)�^��Oj(��y��>@\m�v6O�ɢ�0�UI`��)�J��3�}rͰ��l�-�!W`MJ�n�DW�`h*����z\s�>����o٪�)����S"x~mG�r��y�㿈�0gޯѸ����:�;e������^I�@����ҦlS�
�;��8�8��)�/�5��T bN���f�Ufa4�$�P B0�����uF,������Dn���89��oUj�F!���%h�Z�c��0v��tƼ��<��6bj�޶0:?�F���H
��YzzP��\�{�������e�-\���TT�`�No��ÒcP��!�K����*R[6�6��H3ķg�n gE>϶`+�1D�ë[f�	�}�b%�����j��!AJ�1:4y������|�0j�.ۈG��{��#�$�,c�I%.*��m��# #k%��|Ǟ	OKh5L��� �i���o���ö"od=�ǃ�m�	͔=�$���8_-�����2�N ���4��I�S�;L��w����&�ѷ��H�iO����1�*R�Q��]�z�	>����X��Lf��8	i���i_Ȱ��j�~O{��e	���iº�;�^`��<f��Rtz�܍�}劢���d�C${vNWOST�xXy�3��_x\�b�b��dz#.��F��h��� ��E�\�*��a���/*a�U^{t�d�r�;��SfV�8��G�/s�������
cG��@���8(T���Y@�d�:B�C��kI".�jT�����hiZȧb]�p�� C�.d����k���m�7{�_N�孓�f�8����܀�
�R	[
�[wJ��d�~�t~�1L�9�����8MG�}��x�ڜ�b������4S���1�8�#:G�H�s��-*�e��µ���}ى0�E��P9@kunU�Q�c�D�k<:����R�1���Z�o�'�S|������h�d�Xr]�a?^p��	T�RDgG�$W6S�٫�,$���VL�����qv~Np�ϗ!��b����핰E��jz V�EE��
��a������}6�Z`��d}�����R�j@ui0c���wd=d�1��Fg1�]�*��7�k�딸h%�q�m��耴T!e66��,�i*�ˠ�na�:B�
���Iڪ�<�i�⢓J8�5$����}����	AL�"���"a^��8�Ci�g������=_�.��n��
 �.KL��Ai�gWu����~�<�-�aߙFŰ��'��!��a<.��L8�m%�g�S�ylC�&�����R�`�������q)�_�Ξ1E�nu�.��#ʴR�p^3|��'"O�ޕQ�| K9�
���&UUXQD�y�7�[����<�9��<��,�=�g�86Db�X��"��N"m,� 'g�?y~��޼����gQ!E�^l!7�T�Ѷ��0���%94k��|�j�A�\��?�7�����R�r��!�R�p�#Q&����6����ҁ������ �w�����㹹�tUyU+K���ɸ7�"����:�G��D�[��<\����h�LJ?tli�= �nM��}��O5��]�K38�������6RU*o����H&�!��	23��-�-B�{�W\�d�iK��>1�T�h<��-o	jM��U�Y��B��_Y��D�2Pz��z�$ԁ�[�Sȋ{�� ��m�(n-��p�bu+�E�v�G��G+.��	�T�?���!?�#�u���b��C���m�7�E��WϷT����A�������o$��='B���?nN=|
R��g#Y��f�j�t�=ב���T畦�� 	T��c�P�5r�8�:�,�c^�IƧ<�&h���Ko��������g�a�A݂�&�pJB���a4�(5�=a�h"��5��lw���G�2����FG�7.������W4i�1�W��YV1�$)���%��
�>�Wk?�q���5OS2p^b��9�ǚ����oM��#�">G�<����X+y�R;�~3�����PZSR��K�ApoWª|��������
X7�i����Q%��A�����%2es����Z�Ҹ)��K���N��>�^�U����ED1�`ݿ���Y%������]���4\C���&j�z���Tg<�F��	F�et���wL[ g��*!^�ִ�^��!����X%����i� O�.�퍰�ΆGa�b�#.L�8��i��	̐i���x�	
+F���������Nj�gm�S�6D�)���ځC���� �j�	�	;�`Ng���(I���w�TڋW�Y.g��,Sv����[q����t~E�/zx��6CI 2�9��\�oޑD�����x���
B���Ry���T�|������	�Fr��l�\#��#"l��ږ#����NB�� Y�s��>� ��a��Cg'�O���`їQ��|x��O8ős��oY
�N��� �a��=�@]#s�މ�Uu01�ǖiU!Hea�P;�É����%��!Ђ�$�[��W�\�`�����s�a��7g�F�Mֺⴴ�&��4����w�?F�5Hm�X��0�+�IZ�EN�l8@�Vkf6
������H∼ﵦ��>���9�8��%�� uR�r�ͭ��=.��5�4�2;��O/���+�s�Y'b�ilt���T��l��B�0 ��|K�b�O#,�|���WG��ߩ�M#CG���I'_�j̈�DPXk8vk�(3ƗM[��:.�E!����ҳ� 0>?�8�_o�m�b�������s���v!i���8k ����շ�b����jm���RM�Q0<���uUB4���ܓ�.���M⒛�����o}j�g��]$&��WX:,����?�������7ݗH1VR����{���+�X?�)e��?Vv$���F���<�6ُ2$7%�d�{Lc^�l���R��p��T�a �c��V�E,4�!���q2R�w 2�6��m����]���pJ�\?�Q]`L�������`�$�Y��&"��hL�b"M~���k�@�B��ɥ�]� ����.�z+��F�ƙ���z����)�:���s�ɞ��Kz
�igg�|���2l����/L�)�+�w�7l���K��ٛ�=FF���>n�͝��'� �ag��[v8z�|}Ks;��t)�lxH�X��,}���AY�B����O5yr�*��e���A\���l
�����2�,�O%w��&��3�Y  orAN��LQX;�(���"����/)��55M;s��_��U)[ah����G"�	`���݊dd_2�[�-���}% $��K�#�1Tmu���m��&7�6X��c��.��Ε:mH�/DSD�����T"��7Ă-�2����Ws=Fb_�l8W�>���䳁�ͽ���Zc(�\]�[��-$�b������)1B���6���X�ޭ6���S�sj?�Kg�RP3������Tn?գ~�4���B/�Xa!�۫��2n�e��L?>$����B��b
�~d�Z�T�.{];��͙_�~)0Ld�C7�#8�U���������a�����R��-���S�9�5 �!,�[Ђ�TeF[�������q)���b���|=G !G�`F�	����o�f-G~�(-Oۖ�/�A�/?�O�h�� ސ�Gޜ��b��/����?Qxn�a�T�ޯ
�ԓ�:�$չ0�7di�Ϳ�j�Pϣ?���W�2*�����'T�1���
�w�_sXo�O��y�wXFUY�,^K+�c��^%�?c>��E%]Ok���ɐ﬚uaCb���U��<�઀IU6zy!��1��_�I���	��oؼ�Mҷd�W���mr�f�̒���s��$��r��ߚܫI�:_�����z�="a��l�KkN-g/�#;֝�B$ 4���Gr�f�� m������u1?7�L�����i�uz;E��]�D�o��2ڷ�{����N� y{�nq��ܺ2�ܷ
�Y��P�%�稺�j.�o��%uJr�SO�{��>��ÆS��YU�.�;'z���
yl�E�5��8?�`�,GD#�����fb��A����(�W��t`j�x쁜M
�{;g/��1x�^œ��e�Ab�g��Y/ăގ�@>v�!|忳�1a�(��vHLh���i�EP���b�f{o�~7g��u�]���T٨�ք��~��ڶ��lD�-��qM�}�m�������>�fd��>�Z[��Y����C�N*b��3�8���N�B�zlN�.����ǥN`ڦ�[LN��nj�S�K��B���c�{L�.\I>�D�Ѐ��ʕ+��nb5w����D3#�\Sm�b9�5|&#�*�n:媓�]��9����$*:K�ô��o��>VG��1���q��`��N��H��$���>�׿�27��/�4!���3����	L��q)i�i�>1�8��n��@Yy�mߡ�XѸy�ek
_~�]�6�Ъ&d�����(��9�u8F�#a��O�H\��_yڍW���װ�|�s �b�WMRT�����V�o߂%숋�E?�x�9�y�	�D.[D���[N;�I�,���ϫ����c�� �Ea�(]+$T�?Uڋ�U�c���>5�1t�w�����]�7WX��J%��q)z͇]���!`.�ø�F���+��/��.�v�u'��`�L9���u��I�;<1��<)O!S��8ۧM�PEͿ�o��o���q��h�g��qqT5'`��3z'���}���t�*�v�}��XxB�y�T�0ؙ���=�&����]!�~��&^�黜P��D�o�0Y�#߮�U��9�A�3�ˆڂ�l��e���,!h`l;��\�1c�7�k���:�!��$;�d�',@a=�?��7�V�{�4�m!�/��o(Q;�Gّs��d���`��ЕPQ?�~�8�
������\��W�B��~G�~6�x�������u����^�C,��7���}j��I�v�H1������*��s�w	�G*�ˇ?���quZеm=���;q�ܔt[s�3���9�w�<�^�˹���N���փ�ߒxñ=�n�|E̢���
iuT鑁����U��o⩆UH���xłstzP�ֲ�Ц�#�b���[J|�����w�A��1�Q�R�b��CU��l�v)D�ס�l&�Յ��8�?{jl]X�k徽�S�,Sq��28����V����
�@�ⳤ���:�/��w���������TC�����^���b��W\�)N{�7ْE��=�%�)�{�K���>���#�ܳ��\������f���?�,b6T3��\��k��ˮM>�8�|7%����sT[�I�/���u��_3}ƕ�1|�oL:��)�Xb�:����!�&JI����!%{ǎ<4#��	Cs��c$�v{�����j�!��m�ڭFx��L�t�Jv�@Ɋ�O�v�����s�v��q����y)i��NY��6��Ƕ���Ssmvl�"��#�aAŐ�Ze�vr+�pz)���8������Z
�a�a�_y��	�=� �g��$��V^e3�|��yG�։���r&�z�h�~pY"�o�Y�1�!����H�B��9C���6r+�^e��1�=H�4sX3D��a���hk��>2!㩑�:��h<�rP� <)W)�})�A�;Ia��UI;fz<9s،2���f�� S�l��C�<���_�|;k7�vY��:0��Q��LY��/Җ�j̼�@�	��������#��ff�;,g����&�pN���9-���1�s��G�x����9(�׽�E\ί�j�MEw��i���C��g�W<���������?��)z�%�����i|�)����0t�K�m~9���}ܩ>�ŀ"��i,6���׳��eI�zӂ��\S���_f�E��X_�bğx�R�Pf��֎ ��ٙ`��+���i5�V����h�z���	m�/[�4& �2�U�̧�Z��f{��3�b��*J\|��ȸ-����A4^�>o�U�)?7X>��.�yC`oM������Cem�7!���yF��qFpb�B����j�RdҢ�Dm��8RH��u��up��,���D �<���QW�w����K��=葚W̒������Q�d��`7ݵ�Y�/��E�����(�kb{�z�7op�_� i������'d�� B0�ȫ����)�"U�І-!�.nЯ&`em
�鍈��$�q�{�kc%5��er[�����@C�����X�A3Bڃ��л�,%�닠Ьҟ�����ʱ�;�L�랤�4���l]ݦ�S���~Ȧ��"���0�H��s� �tD6)�$�#q9j�����"�hBi_8�:��Zb`�'?C˪�Y�<�'����zD_��Ѕ�$���Z�O
D$+�P�c{Ў5:BI �7����l���ծw�%N�68l���ZI˗ٖ ���6t����U�*/ �h���?m�eG�(E�y�0����O\'�����0.�z��fNR��q�>Ձ���������䳳�y���D��Y���s�Rw
v}�����d��:�:�Ex�<�V�!W��]��̞�� y:OJ��2��+��^.k���Q�W@��%b�*l�H��2N�8f�'��u|: "����.�D���ȕ�2^k���I�/QԻ��X�q���im[@���ؖ�8����v%�[+>˪�2CO�!�$w���ٲ�Y�K��*.��;5�c|+�=�1�x~A��Y�+@X� 0H�$���JM�^`�Xe9(J���Jp��8*;w2�%����]� $�P��П�ds�䂟�^^�n�E���6����� b�F��{�dڷ��z!���a=(�%"��.\�ؙ�P����׌v��mP�R�ɸ����-�Z`�A��y$) T�<}��z�3��������kzN��e�Ͽ��Ȭ������Yt�W!o��$/zaG�����L�ϭ����1ώ��ee}��}	 ��O�n�>R	�G>z�Ճ�X�v�S�k� �:��'��T0a�'5<���y�a��ih$��ȷ_��JxT��#ƏNˍ�_Y��1%��f�;�ϊ��Ż�Bÿ�`T�p�3�1~5�KПJ�oY��l�ס���_C��*K�D�<�W��Px���S��Y���(q�x�L���U�F�c������5�������z����N:̊!Mb���� Q4�Hz�Rz$���VV�R)_����նF���ҢA�-�-�g����������b�J��<=k�kT������R�j��n%	p"�J�-���ڲ �:֭�{&@�f���ꮋ��N����4v.��ZN� y����y�[&��_Zw�D<\v;כ�Ȗ� xi�z*�a%����'Db��ߞ!l�W�W����Vw�� ���:�凮�ӊ�����~�̐]
�T��9.���i���Rr�^ ����'����!D^�@G./1�� س7���טZ��J����#͕hȗ�(�V����?q�K��R).�������>	mc�p\�B�Dsg`�(�tP����xl�����!�F�gǧ��'z���n�Ծͧ��}zDp�����`��]�H�",�Do�f�~��<��2����@�1�_��Yso���}5���qISvA�l�[�m�D�b� ��,�����z_f/�Hd]%w�<rQw��W��烜��	lB����"����_5�O��"	��RB#�y��
X#��� ߐ��R5!;Ԑ���	�ٺ�ᵯ}�������d[�����׾qā߈�jn��i��\��"rrc���14��c������x�y#Gɘ��"U����t)-�$��Lӹ����?��1Y�D�S<��C������#��~�}U�hr�r��;,x_4Rx@V�Af��1`��	D3���.����m,���Ѝf.�*��[8�N��@�"mm��y�I�&��<lG���<F��A��N3b��p�K)�*��=��2� �2�H��@PF=�W�Tt�� e\����� A�?S�?�p�t)�.�&3ġ�m���^ɫ��x%�O=A�A\��پ	�X��F-H�iy���g�{6��Fv�EŚ8)���'
0)Y-���M�r��I+=A���հ��Z��9Rݕ���9�?ZP��kr%��^3�q�S���]���5�ɽ�<�y7D�[��M�v�*E$�^�z.�DY��V�3��n&�eΣP華SDN�	)����63�%��w�@�<sU+�I����dn�eԾ���M��b+9=#�����C��Q�`����v�J����sM���hP��Ҹ��~�v�{�N��dY�]Rg�Ȑ����Љ�l��V��>>#�2�]%���Ce�ߙn^UE��'#�u%ϳ͘�wԁ�A��8h0뉼��\�<O��$�_$LA���NQ�+��P����"�ڇm_Ki������GgL��'��t
	�I�}�bH~ﹾʧ2�JL���Hi���f�%m�g��܃�6t�dIj��"+�;��vgl$G.M i��`���v�v�^JzH�e�������կuR�cw@���e&���b²��p�/��I�=��C}�@��O:Z
�������V�=_���K߶������ �t@{	0���k�L��3M��5�`LoJ^��2i2���CU��x��޳ӟ��_�ф����3_�Q��؊'���2���E�S��eT=�l
C�N�Gƿa\�W#����<��[�xr[���:LE
���IJ a�i������:�%�?>�7�^�Z��B�vS�k�/����q*�L����U�rTD�r~;��#��ӧ�����!�N��*Cp	d(��~��[��QwrY#K�n6\�z�y�uʬ�B��u}��p����%S�2��E،W���H7I���Ρ�2�m���N�fv
t�0����5[>��6'�E%x�{���,��ͫI�^��L�煊��5�T���^p�)�R�VD9��#56�P�^�:�K=��TTO��D�pݬ��%�KQ��O�0�q	9�P�j�J
8��[	�����u���'��Dǡ����!�,�AuOU�Ơf��ۆ�D����HZ�N5Z���݂�_e/2nPU҆����&���h�ܙ0�꺙��K���B����>�#綣x�,��5h�Q'�ŗ�ᕈ�g����~͈�6����J�,y��(�S���ڔ72E�OdΛ��r�}�m����|��E�z��m淐�Jzw��>ϣ�{X�?&B1Ӓ�)�/�'?T񪅐��=cG�BkR����PX����sS1]4t�]cC�TY\�RmH_,�c �'�LN�'����w�^�kU���ڦ2����>b
1����+�|�V�6iN_A\�l��ҋ1�=��=��:��ȮQL��e����_n��{��B��3���O�KPT������ P�����)�6�\Vx�e��o�Z����8��k����"+|��/5b5���x���{�J3v|�ve���Z^;T#�'��T@gK��Oy~�s�'�>�q��mפ�����Jrv>���d ~��[r��J�_��迢�z/���FL؟�v��Gز�\j�S/g�_�H�+|���K�"<�}�d�y�e�h�t��$6�:��^�7�iS0]j��pQb��z#�)��YQ�0���}?��aEc�.��\hT�%��G���ʨKF��%E���P�O�:����N`�@5ې��u �4�G���^����l�	u������v�ٚ/��Du&��=�����uQ|Eey�P����#mSca���9��	ſ��b�t�͚)�{pMY�����ψG������m�s8Ȃ�љ�ʷ�,��%{.U<�� '��5��q���̐*±"��%����u�b���}$�+����uM�ne5#ZO���&���ji��<3D(G*����j�����fu*��Xsti����|(2��F�C{�l^y̲�??Ui�()
Vhh)]���M?�t⧆�%�в�1��?#��r�tI��Or/G+WQ�:0�����5U�;0/���Q�v����ػ�x�p#vX��x%ҵ��o01z�aj���[/1�P"�<?��8m�6YO �b�n�:24ڡ4:�jݒ#y/�]��4-�Ƨ�ZI�}}�FWc�돦�]T���>�g4�(u�"�����[�EU ڲ�+{hx�`�[F��} 1=<���Ct(�����_A��ǆ���bd����܋Ĉ?q�"�����G"�9U�,:��D����#8k2�@������[8�o#�'>����zm����4Oha���gi��n4G��~V�s��O����]�IC�cĢ�-cy]�]h]Vr>��TjT�L��ƒ,�Jv>B��h�&�.V�^)��tE�U�W�uL�s?^|�S��r��K�J"=TR����p����U{� 3+ގIQ��e��<͐�+5|�8
��B��)U��n���Ē��[� �2�G޼@��]^4��A�+�9�=	�����W�Ů ����F��l<��ʃ5ó�ʠ���d�w֌��-"h!��~(\S���5���dLh{w/�&�V���ɿp���#{"�*�+�E{�1q�'	�n aT���^����1[HhZ0�K���{��U��|9�V��zL|��𥵮Q@K(YY� W[W[�ò��rb��h��j�I}�rްer7�G%�_Ԉ|�:��Kx��r�8۪+XV� =��0*���K.A4�^{B��~{z���Pڂ���JU'!|phgF�<yA�;�`Y+�Y�b���S�I�_KӀ
�t���*{������4psj��N��!dJq�Pw�[��3�X2��~Bj�Y�����Ed*�v1�`�Ji�UO�(����^���vc���.�+�j1�{���j��\v�W�@����*���tG!E�}I�����B�^S��'}R7q�ޤ~��3�6�Jм[t��M�ѱ>���^�`��:ښ
��\X�R3�X.s ���1#�׋�����g_ҍ/�F��_��OZT� >���������\���j�o��8l%_�Sԥev#C��u7�P&`�-�;|-�o����N�6�dl��D��hC�&|4՟����?��s�ܱVL�$�rP	|���(T ���Wi�+L��mB
�&��94W*(�����[ﾫ�3I4��Ř`)B�U��uW�q~�6�+���}�)��N��b�u���ĩ���z��=0�`8��� 6VOF�"�C�ƻXC'��&"�u��?"��{���ǥ�"��R|m)rؐ[z�3�U	�ȩ�/�+x��P�43��Ƞm��&N�TTa�qk8���P)�Ze��w���v]O�`��B�m�)9ѩG1��a�͌$�С٠�wA8w������|]����\�\w��,���S� �g�w�h컵}$�JI�O|�Q�'-�
�ҦT�բ%�$Dް6�>=�5���ڙ��� R��e���� $z*��Rt&��WudW"�DQ&��Uu��2*1�_V���2tCG��`|߳˳�߷gtS��t8SO��OnR��&�`���R��K�/$��U�CpV.��S�b��*����B��H��PΌIl��ՓY�2?���� �o����m��ex3ז=/O)Ъx� �*MP-݂Q8���yf{�D��X$]�m2��(~:��1|$�7�������Q�zx�U^~��R�Gf�eb~�֜�1�{c���$e�_:(I�n�D7w�{��`##U���8�P���X�m��#�&���Y5�T%cq*Ϩ���}e����#ß�D��|$*����(V�j�H�w��0�X{�B�cD����'��ئv��ʥX��O3g}s3ÜR>���� }t�7U�Q��K��"����`8��h�)�s�2�׋f��Q����)��W��v����M]e���y��G���iXB�a�O��&�����`�6w�jW�H�s��#��'D��&���V�Y�W�����iL@&U�tg�x�]|sz+��Ꞔ n���/8#���"���OF��,��g�j�B(8N�&sVļ��M��t�=��l1eM��i�ߪrA��t�����xKQ�Ic^�	A��R���y����_�pࢲn)	���<uI�]�לL� ���|6��K m `Sgrƶ���l6��r��&��`-�`\23*d�Ǝ$�4);9� ûF,��ȑ��@�i K�Ə�?����(��Y���1�����'\��An��v��qh��� X[��t�Ո'A�a��*�UH�o}�n�m��X��	_kO�T*���kKdEJ�x{��5\�)X�l 1�癘a�ݔ_��R8[F�n� &��:h�Q>�ן���?�_WF2Bd6J��.�����:�~P	8����c�c0����!{�UD���'YQ�fq�;�Vr	8����jvd[K9{{�Zj��&�ug����j�<
�E�|qǂ�X�ɘ���:���i���_�� 2��5pHə�<�r�U3q�D����c믲��~A��!�DĂ��ե��y���E3���[�޸��Rk?����L���4�M�t�C�J��N�/И�((Q��bi�<kr��c!����lMmE"����q����ْ=%;��7n�DP��ɬ]jŅ�CC��Û��è���AW-�wt��$�J|�dɜ��~fxm���*��CbC:b�TS��W+!q�=/u���Z��:�h#���<�KК�4&b3z(�v(̭	zu���XTZE4��|� |m�c�s���>�;���c��6��AR{�\
`�xt����B��P�����s�RJ'���I�[�B8u$��g��#�c��t�Gx�g�;,�}�Evp8��8�t$�G���~��d)����#��@��խ��f��* ��[Ε�������*��U��a�c\~n��ښ�v<�_�>��{�OD�i3l�Ը�����-�'7q���U=�;uZ���ʁ�2��`>�/����^;R9/M���N���(�d� ń�+�\S�Ts���@�5]���!�S3��7{�"���z7�6�6T
ݡuO|81ܤ"����m&���,;�;n厜��,��;D�d�no,	�3�\�#_�أt6��6�}f���+&¢����W��b�x�֢G� �4�ؒ����'����9����Ē�xـ'�X�PH�rH��<�u�Fw�e���K��� �''���;�ٕ3����W���5�=��˾�G��1�
<�x�^1��v���A��ʃ�ȹ���Dt���2���5�c&2f�6���z��u��i;@�	�<#�M�٠�r6l+=Mz���	hT�r��l�qC���|$!�W�=�_4���?~�5(�i�9������]�@��B��.�^�k�� ��X1��dt�Q��[˔p�z-��j"�O�nR��.4��t�םPh���R�K=rN�U����P-~��xKL���1Z�,�Dr8�`�,�@g`���;~~� �GΡ�%�+�͡��n�+ᬃ앸���c@u�V����������ӭ:���&��l�.&�v}�2�w���۷�x�
��7�c>��c�_���������R�9[���[ְ�,!~��0a�K�Y$:��1L��Ϧ�B5�*��5N��<�����0������e߱�e� 3D����������%ŋ�3�b�w�r���|�=!��|~�E��BQ �"B��ZT��B���cUR s>B�ϯh�"�7pT���ڊ���u�HL��^g��5ئŅ��9��Ʊn3"C�<����7�b
8>��ĉM�<Y 2��NQ��^�����T:�j�K�U*��'(��FM��zz2xD����d��� r!�3�ձ0�>#��Nژ7*hІ�<mG�`1N>�ӝʖ�����-�ݐ	wwEiU)E��ڛp���&Pd��㜬@\2;�JB �u���RFT�SsǢ��Sb����z�%��Vvn��(�5�<B�RŁ
To�|!Eԧ�33����=7p��W�[0q{�yUrk�)s@H�l��[�L���hS1����ƛ쌩x�x� `��=ò�5kL�jo:��?���F�]�y~��n\�u���6Bj��Hn��G\fK�S2�x��z-������1��I��C��G(%��&b�>���b>���w(mڿ��Z�q�ٌb�&﹣�0��9�fخf�_9$L�}Q���Pɻ�}j;Y�#]�A{�vA��X?� �(����P�K�\�Ӛ�<��5Pƙ�uɈ�(�n�����R��#�����ͦ���kP���(�Tw����zb~i:��9�f�.>Ls��՞t1u+�RYy���=���h�`8�ee��{��-��V�K1�3�v�W��x���M��YR�M�t_J0:R|���~�Ǥm�E�	du��٠Nz)��t��K~jl�OY3�;~=�w�`���x�@r#}�+�N.^T<h��ĶN�?/��k�A�	L����`6��N?ۏ���苻JJ�(��o\,ۇ��~�����Z�b
ՠy+L��JgH5�o���5HzG���~���`�H4�d>Fgn��G��p�&�6�0�4��E���&H�4����U�TՉ����ݺh�/d��-e�[/��,��J�\UHz�KM(�y(�>i�W˔M�Q�
v�-�ˣ�c5��wT��ZU.��[-��_=���%�+(s��U>�[�ڒj�ׁ_1~q��r}�D��A׫˼�;���هhxאҝ"(��lOR�~~!�?-�xF�@�)�\%� �J�Ѭ�x<�����ـ�l��s��y�:����+���Z�|�gg67���O 3���y�au Ʒ޵�x�¹ŋ���;wҪ��p�+���Ip��6��Ol+�o�WDH���cW�~vUO;�O��g~[���� �Y��N,Y��k�M�v��1�[%��d����o*�3�>4����d��$T��\�Ek��.�'��Xu��uAZ!��B��$��I�~���vT��U�x�{ 2�˕������?�F��(8q#<`��P�9-��l��t�S#�Tbv',Jђ�*X/;Osqu��W��W�ˡ_�Ϙ��dK&�Qd�}��L
��6����?�2T���:>���?��n�&�GI�W8lv�9���*�m=�\�������q��U��q����>q�կ��tIlk�Ƅ��lg�b����TG� �����m�RY�X�w����E���7�b��O�����V���flI�E1v�q�7�s?��V���R�/���V�>��w0A�u�5�/ �g��� :��@��f|�觰T��<ʴ��g⼷O�/��c8���*�9��:��+l�,[��+�������6�E�b#�(���I@G�?e���޾��~�to*g	��tG�������&B��dK�B�yT;�_
�FD�5j���2�r�� �-0�{`�>��w!��"�waPmI���JG�6���¨O�'j"����ϻ����j�6�YK��%H,W.&�8Ҷ�gѷ�k(����aj�KCo��,�d`�J�o�3���M�����lB����R�����n�{��;����B��0ѕTӎ�6�Y�k�z$y�#������d���vL��MJ��jg�<+\I����l8�J�`�OOx;ٮ�^n;�0�4�ӠXT�~U�z�'�5������'�. a'8�p;c�~�N�et���K�ei�tD�D�%k4.�?��p��5�W�П���Y6�'����7G�����TSV��Q���32�pSI����B
����Sq��t:�-B������ѡ��궈y^]����푍9�L�4�
�I%*�@��_���4�T���G�A^�Y&]�޿�s2���}WT�&������#?yl�������M&�����U����^�<ۂ���k�~�$@�"��~��ޱ?s;�*6���Z'hR��S����u��z߬���'��(��@6��m��|=�K��*��"�5@:7��-=���֊� �\��ܽ��9������6%G!K�vDV��EY�owt�ٮ�#O�d 9��S$�^0��Rۣ��8��'5�k�b[[_�KD����氒�Yb�|Ԡ(�ҦW�0���meO��gO���A4�Q����|�_SR�|����ϡ4��D�uyL2)�ǖ��@�{
�S ")I�]Pl �#�~��0�`K-+�N'S>�]E�||Bq�����N	�)A�ͅ�_��E���&�;�w翄^��4z�����(R}�y��\
�Uj�$���Mh�:�|г��L"xq30eBm/u��g���q��/��
{A�c�S]�}��/'���&B�*fB���Մ�4@g��ңn*�d�����ϊ�`��W8iـ�Y�C�[�,OcQ�>����>����|�� �K���N�� �J;.]��;tZM�i�Z-- �F)��2����L?_�9X�0�c7_�(?��D��ѓ���+���t���p[&򖣙�y#I6�I�j_,�W����&~������b�c%])���.�7>Q+%O�k�  e��H/_��M]�qۢFXN�ޓ��������WU�˔tc&Y+���,��\2�I�m �����0YJ��Ztb��׵�2rIDj��S�ߪnz���Y�TM�(q�P��+����� ~Y�[O���"�\��Ki�h��d?}&�(����b���K��^��nAGHۖ*�B�Nܕf$���X]��*/l{��E�����_�m��Y�bΏ41�ojν�]����l<���k�l� 5ȟq�U�o��ϠK�>����|�z�t"H{�Zٙ��>���.�;J��Z�B6��LϨ�Ur�"�C�`���"c����9a����g'�.,���p��#�?�����0->�P8�*��9�:V'�|ny B�L���#Hq�҃��'1���L~�x�u�P��dU"�Ȉ�w�N&!�>ŀ��/�Z�8t��m�k�GԷ�N�	l�� ��S�.B��ϱ�u��5�\@�����{�?_(=� �R�j2{��ڎe��oϨ�@�q�<1|�d��<������x�'��Ƕ�^�GA�ʒ��)�4g��
�_�]~�ŝ�i�pU���.d����4���>y�0���cL��x����R��P�:֪��*a $��˷G��D0��l㐑��E(�e�{,ԲEX����z��2&]���%� �b�5�Lo/xݐdB�O�����t�y��@��4�D��ҮAN�
s����#5�8�)F��j*�:��6.jv����#�HAҪҿ��}|��(G�q8> s�.t|��6@3.H|.�zm���3 8h�a"���?�йV ��=�Ĭ j%!=N�t��tS����%x4h�6��h��.�S�Yr���M�ꑰLS��w�#m=���0*�qM֡����@��*(��em�<դP-J�Q q��׽(��0�ׂ)�ސi����� C���d��䥕qų�������!���b��:<.띍y�b�@XH��,�[}����N6�Y0��d���X{����ZB��]����B���E�FH����b�N.4h@�`��Rh:��~6�!��¤30%�t���y��C�@Ͻ��A�g�ۼ|>�Eu�OџpNdRP�oW��ei�%�B�`>������<r ��P��&���}���X�8��9[�8�g�яf�Cd(��{�H���u��vIC�{��K�'��_�O��M�I��x�Q^2S̥0Z��V���	Yz���������t]�د*I�h�C��Mh�v��X�-a�x(���Ⓐ ;V�?��Y�Oa�k\�ա��s�P1�Z��{��<3`�F���b't�<�`�7��Homvw=R�6�.̆����ަ����[��P��|�2����y��Չ�30���i~��ҞC�.�U�O�"��O|GɌi���5|��@��/��J�X�+���Z�Ejl_��ۜ����sT�R�[�n����0�M:�����κ�e�Q��P�y4_幪u�^�d��r���ј6�>�u�!��f�H��t>b��Br�9Vz0�P@�E���&�5����I�%�r�@j����߭V2�O4��w�Aڟo�LU��N!K��آ��6^��T�w2�>k�@����"t�� 8s����xR��{�ks�ߓ�\��Vt����H�+K����@+��UsY��-Y��BWX�Mq�^E���?@��m�榝?؂�~�֡�%D�S4r�H�x4��^+��^C��L�9��?������C�40z�e�'�ʸw�'��J��1��mKk�ݛ�MDJ��=_�����rӈ�3�6�8[ YX��>O�τ�x���eD:�Cl�x����X�������N�6��?��=�e�^�/�bL=#���^�������bD.X8��@b��A��H����SDm�%��J�U�"!$�n'��,d�נ�Z+��&-��p`��M
=�o�a"�"�㟫/�!�ܠj�.C��P���T��/�!b��ta��k�<5H)b���Y�D9��r����&��z��z�z�@!C����$Bw�F^X�щ 4>�(�����0a�9�Do{eN��]�'���LHn��f?@����,����*�\�G�ٝ�4k0�"Hc���������s�`ς�L��uSU͞�wkO �;� 4�+�N��3����ެ.��1Fk	�o8"� \��!�Q}����E.R����Et���XU��>0c�@GfB�����($�����+s�v��d0����C 4�<�����P�K�U�ò��4�b�PP&[q�5Z�
��v���&]�?�gݩ���c�
���mO������2��|�l*jL�T���@��Փe.Gかy��\��``���I�0�u4�u#�j*��f���P�=U7$�Tj�2�jQ퇤����B���~bD��y$�C�g[n��˷�	��XDfӘ?�5йg��,�??;��`��O�-gpW��S+.�4ح]���?0�~Vc�m�������}S��øra�fF"�z�H���w���Ǌ��Ք�����c��t�Bu��x�4V��h��s�!�fp���_�9�YFY�� ��ĺ��u����*S���H8Rc�4xQ�D��?Ht+^j�u2���Qc�z���jW���(\��"���-�tj���q���>Mr�4�|3S��N%���������2&u%[�U�bB�ˡ�HǢl�ӯ�y�@�J�9)bv��닡��ƽR�܌��A&��Jۖ-��+Hm�6q��y���l���5l�bq�A��u�Z^S�$�
s��
e����U�2롪�sV|��	v����|��1�s(7�u��~�FK|=��ڳ�8��<~N�z�؆KW��[��c���M~��}ޞw�`����YN�����\JZ��j�Eo���ǚL\���x���M�{d��Tvvk�/Ǩ^�'�b��+�k��F��KE5]�--���*		�/�a T�%��>]�9a��@֟w�Cd�[qsD?�]{����N=����b�G�G�ʀ�ׅ�u�n�����W˺��b	[7In�̓C��웋2; XL0'���r����@I��3�{s�r8ŵwu�ͱ�V{3��?�[�a�zJ��J��`� n(:��LB���Xɘg��%��I��q�!�F�����?y��L���d,j���}BM����MŤ�tq3�W��F!��Vԕ!�rN�D�vW�%�Yt�����aM��e��@i�ף��0�E�������p~�]js�ڣuלv�`�	�ĥ�X���z07��m�_?VC����[Ѝ��5�������P��^�Wo���ڽ@`���;.�����8��彄ct��s�d4:�$��%*�YS�W�@��z���>��&��0�Ƞ6,�ڦ�f�x0�14�����i��+���%O�
ܵ�"R�\�ed�C�tHt���[t���¢#}bh|��5��`S#NOt7�
V"�;5�� 2���nR����V��(�N7v��"0��*�G��@%>UMg����e����l�>��	eK�݋�0�\��l��U��y���7��(bY���Q��h�л���H'?%�Z�n-0[#;'=��UXfnz�Q��U}~�oZ�q��Q�"�%,$h|U��j*i�S�[�4}��]�}�1�����7�M����Z�Ä2{B}rHZۆ�O{��& ��T"���-�(��6$�l�������ధ{6
r5�����\��u�	u7睪-����-��XW� O��'@����X���s����.�R��0�y/�������h�n+y�����Ţ�e��p�0����4���J�6����(���U8��p_�����0�c^��ds�����0a�|gѽ��b����Q�TEH�tLw���|C�,��&xWu^��vߝ�_��0���}���U?��˹D��Sڔ�8>�y�۔?ň�e9�����l;�4r$�|�J:W{j�˱�<�D0s����u�J�����A�>@�M�x=�������x0���&�z�s��~� ������=Z������:�Y��%�.�͚|)�!_�Wa�zM�l��.`�\xS4$��N�%�m8��!��%�QW9?nY�*±0���m�U��ef��AYIMj$�P֮���C�8O(a�	��+��FM�t6J��v��TbLe�7Z$G����y�;]U)�Q���'�cohy��\�<0�+�|l�H�i�v`1��`�ڹ�{6ҭ��gkZz�[G.0������&��)��ӥ[�4���E���It��@��Q���N�P�ӂ3��8�ۊӾ녁�X�7/	�V�|��Ui��\p������ύ��YB�N@����ӑ�2�Vn�F��nL{ݱU�fM���-n�v��踅�Eٞ<)�7�崣��(�^jJ�c��g��L�3�ż�����p�� ��l�� &��@K؜�Ɛ�s��8�W�^D���i_(�g��3.��c�ԇv�bU��[e�}��r����6
��;�vOiZ��ƴ�j2�АM$L���Ւ��,����������d��F~��baզ<`�F�&�N&�g��6��Q���;r�dg������ #�n��d��EIMgE�_:�(��Fw��U��}�����	�l��&�8�sl����0��m�cu !IHx%{�uP�V�pN���}{�P8Δ�.��mw	�e��H9��b�_��䵵�i��k;Ƭ�gֿ��;���T��/�Ҁ�]���9�%�x��-L�X�k�ԡ���Q��_��#^������
�0="�P�� 5���	�T���1p)�ipc?�>��Q02��m����Λ�H9��0aT!e��J���N��B��B&�g�X���w#X�&~��e�{�;�'�N(#iCY�
S ~2Q}W��#�cl"9�"��p#�'��䰓(��P�s��xSr�(N`����NH!d4�:G�����6&�� *#v���f��3U��ʫ�u�#tU��_:���j|��Mѩ�,	E�������?=�ސYFʣ�j �"
S�́ʑ�_�c�~+�QwY��kg �a��͈�K/~E<}�!h�4'r-<���Åac�
�|8�Er�5No���7ERg�+S��3�@�}n�� ������/����A�/m?��UCn�.�9�)q�>ui�{\�|9��UŎ�kM9��S;��J�G34�e�نK*^A�&&�K����>��1�e���#9I��;������L4�)G�>���|UU����O0צ�ʫ vU��+� �ɓ�{�J�� }�����.���B%�b�=�w�
�����;0i� �[E�L]���k����6u�[RB���!�X��n���R!"��?>x����o���'iL�a6	�?��-ᗠI��C�$>|[]cb1F��_)33��d��rn�3j�1~���k��
h����SȻN�4�`� Y�p��$	$��)A&m�7zUS�9_Ub��I���-+�/��(P�H^�8�<���6 �|v��6b�<0 �o(�]L�<A�ÝMv�";OYek���j��R@��>�h��4=H
��B�vhR�́,C�Ck��]Q�n����ar�o(_����$�ת����NHot���'�'�%3b\	畉�J�8P[�6̻"B�i��iձ�3j1��SSt.T��.�e�IсK
�X�Y���a�FM����FȎ6�Q>L��U:���#!�������C�-:�""���a{��eq�9]�s?��H��ʞ��ᵊ~:��u��l_n�h'��!���<E���U9D�PehXً	�_s�"7@6���9@�Qe,�@��f�[�[�X�&!��M�K����ACvҸr��N.'tK�y�q�T ��ܷh��>51�X����dXH��h�p�i�x{3rb)�Dh���wx��+t�c�G�� hl�!*8�R[N���=�}{��,�g4� ���%L�a5�8Gi�����CO��	ي�����Z��/H�}��� {$��������:�A�[}5+/QSo��&KUn��V�?�����Z�[1��RG�Z-u~:0�9���д�n���-Ɔ\Y�`l�<�j��D�r��I%��3p����"��	�`���Y�I��*�����	*Ȇ�Ùđ��BIҌ�l�-����B�/y��XO�u�xdr[�9����ë� �s�����N�$4��V��&J>� ��R�����ފ���Ў"��႟^��\�%��ᬏ_f��x�F���:��݄��ghG��Ep��K���d0�T܅!��52� ��/`�붦�>����4h���aC�����ZgWkY������ߝ��%��5�[Ho�����d��"�OxWmL)�G�U3~�������r�JЂ�6�J���OU��d"L�nع}�пI��z<Y�T7�/ڣ/�[��.kr5�����=��4_�I����c~k�G�%�e���<B���kNa�Z�R�S2&�5/�y^��x��E��B	�p��"�� j�+2�_�u�^��m���⪾���MDFuH�����?7C��h����Q[ʟ](�H�>�O�����~��װ�,O�E��l��;��%�8���Z�'�����M=�����?,�Sc����֡\	��(������� 4�P:���BN���0�wc!'blq��l����~ŀ�� ��:��A��g|K��N^e���n$eC�5�{\`�#Ͱ���y)F����	�|4�>o_6]mH�B��۳�`�yۄ~�x�ᘰδ��<�+���J[C����.]�ŭO�p�
Vq&z������a�$�s�����e5Z�O)�p�I]�"}�c�뒿<���ɚt_�������i��$��ukB�[@�c^z�(yr,��a��{�?�@+ii)�.t����Ŧ�k���-�Ek�5�-ZV��������7���3�<����e��,�,�$WU�wi�\,!��>5�;sB",d��NW�@N.��ZY����63�߅(r�9�']�XO^�"�*F6���N�PkÉ�W��w�sv�;�E9M�J�ln�؊��q݉�EJ��q��C��2�Cs��d�~�:�+�ڨ��kat���9"�.�����T��qШ�kVe0�&-����)�j�f\�<��5�bj�(�4�%����8j�㝸O?}���$��jpp'��A��8uϳ]�)��7m���~��y�a�R����ݻ6?"��u����)��|o:6�U�bEoz�^qҚ/M$�kź���ؓ+�_���7��΋ՠ+z)�yB��L�a�kx�Q�u��1�Lۿ��2������>R�.[4VqN�[:��C�ON;���2�]�>fv�,���4�=���+�1��Z�PJ����C��Q�s�����
ˮظ��=�3��KC$ˇ�w��� U�$@�䳼��Ma�TڿQh�XZO4X��������s��?V`_z�*��N�#Bd��q^��O���i%���=`��F]��X�{��?[�0��Q�D�Vh7�0ԥ��a�IV�͟����;�̵Y����m ��N"�d ��>��I�QxM�O���i��ۦ�)c�z���E˛,g��r����� ֒���G98e�.X�e��fj����[�,��?�)i���⯜��n2�24F 	7��F(���g�~p� �f�ṓ�M��C��}S�L��|�1T~�c��6��>��Y.>a�12M�Ǡ�Mv./�lX��P�����gt�D�l��`>|4WA鹹�/
r![�%İY���}�d�qב�z���d��5}�W�bi3���6.��ۮ��o#0�\�zg'ͣ�O�S6yd�Xl0�N���t� ��Z1O��#�ݩfV��6�5D�]��ʔ۠��v�R�m��E��C���E�B��1ΐ��j@(��d^�X�����ӽ��Fї��~/1�Q�fб��ޕ7�͘b���Q|O7S��}!q�j=^J1�]���r�1�~�X�I�U)ܓ����-S�C-��c��joe��ڜ<f$���ڮ��g5�ȍV�H��#v�1���^E7S��1��:��|�07�U�[��ZO�׵*BfD�Օs��?:�i���faeJb�o��/s1�E�)�~R�j߻d�F�e�Ć�C�����NX�@�fy=��̳b���۵1JH�b�%�tF�'i`Ѵ����{����u�X�Y�?�%��*QM��Π��k�vK����_��W�gA2��Jc=^w�/���h]֒QzAϛ��%CL֧���@��=��w20���~zY=��[P8��z� �ê\�%rpo���'+]���iyR���9[
�@�����)�7{���;���� �Ю�ҙ�HZ#�ߨ 6��MT�'�Ԉ�1��ʗ����Y�ub�F_�������Bӿ9�����oLc��7�6m�i�~�F�W+��f�z��ƕsG����ZC��N���t���Tm�.�8���a1�0ۦ%�:�۱y$�3��NQ��3ۧ��&d.�ݏv�UEi g�������4�N���m�,��A�5yR��fUP�_\��	�(�ֺV��f��*��^/Exقr�WKi��	���<q��5}L���l��t�9Ĩ��ڡ���%� g�F�B �r���u�e�
�3��nz:X3"��'�|�����m��[���a ��Ԗ�,���@��V���V�N�D��--+���<��Pey���m�1�N���*�^/SQh$�n��.o�1 � ��t�j�}��ߠ4��3�zD��I��D�`�̔�b(�� 8X�m�eYǮh�h���w�4㝶R�8��ę6�e/��[W�k%q���B�������b��@� Ɗ}�6�X�<��?�VQ�;��&p�hC+hH���G�O.-GO���h�/�G���A�R�N������3���ڳ� ���X0�P����`��7f,�!�_�eY��#�:X�`IM���RM�9�g�#���%� �0x.\��c<�'��@1�m�\��E��(vk���n��-Ƥ��OQ����5#��$����C�a )n��}�M�jYn�8��ْ�?(�{B�#�)z][G	�:�����N9*rS��T�t�]R\<�#�u�R*��O]��N*5MC2���7e��m�7[.�����U,�ˏ�a%��U����<}�S��og%}#,�j%�f��U��<��p�������>F|���{�F�2��Ę�Q�R�t'���*���+��veGc���k�(�����h��)��M���"��,}���i5B*0.��l��% ��S.���ԯ+�������.����`ON��F�目b�%�l;�K�9)�?�w�'�h�_5��I�tA�TI�t������k�/��Ě���b�Θ��"�ɽ�;�����o�`2r�V�#s�%�Wh����ɩQ{�$A�6 �6ED��H�jms"=���dz�Z(F}F�卻����66�����߻����W�Y���2�M���`�跡x����+\�E��R,H2��rz��)'�Yf�4���z?�r�����S�����hv��7����t+i����Z��W�w&`Ax+d�93>~t�X�ūu׵*IC�W�OL:��%��@��)��"�|���Gu�8���/��4�gt�^q/NO�:�V �6�f�$RQ�χ��-ː���Wý�N��TC^7���q�KZs�վ��Z�3n���Ծ�<��r����ICr��+�׎(W3��`&O
q����H����$o�o�4{լp�L��Dn��?C~.�d(ٔ�'>5s����*;��9u�Dt���T�*-u|��1^�C��Z=c���,��P��%.Z������,< ۄ%�Ģ�����CغD�}˅3mx�p(`�������cZ�*uw�΅O�Q�>��H�2�7\�
��/�5��lո�G��'�m�D�x���5[OKw �y�����g��� !����Z�8d�*#3-+R�xk$��Z/2]8¢�"N ��7�!�����q�p��M���o�BH���k*���9��L�/T8��Lz���r��97)��(+}@����"�3����K[�I^���i����@u������%�k�iI�v�&rj�aBpH���i�l���6&-F#4M�Ae[O
�BIK��tf/RW��;������܎�������<֟��Mۘ3������!M��^�����&j^|[��wg���f�zp��'�󪜜�D�N{�/ϸ�8�-��D�#7�]��'�6�+[������2?MT���Uv~:	U%HxEH�ߙ��H�_��[@��,��K"��8YO��D�߼@&�ax�F��	�����9�)h'�*F��[	J�<�u����D6�]J�������Ub��(�*�Pp6�uGx����,c���yKpc��Ǭ��d�9��#M�o�V
�VT�ٗ�%v�FRhe]!X��/��H���K�G4����#Iu4U�*���r8ˣ�� ��3/@�κå1:n#G���4�2�Lm�ݖ�y1����H�����{D��_��W���H�wi�2(]���m�>7�_L�[2K%����{�L��Y3���yr]5��Ux�c��a?D ����b�1���Ÿ�LF�8��<2��dԾӻ���l�sv�u��U͏�1��w�+�sm8�1鯹/1��Q+��/��ʘ���
���8`�����«3>���S��W��W��*�%�c�\C QG~�c�;o�:��{1oC��GLO�
���Ñf��T��\^YP��Z��E�\�6rK�N�	�$������X����0�w`=|��E��<w�X���ŭoJzVS`�V-�	'�[at� ����i֤�Y�#��.���a
�d�h�}�&�X���.8	�����k̕����?��n�K�w��Y �Y�x~g�d*d!��Þ��~eU��O�W�~s����Gt;�����LL�3��NI��#Z�%K&*���\���(s�щ8b.V�T����3�7������X4:�׾�������P��DH�F���G#�k�WË�Ѻp��z�lNm�&mS6��83�)���A%�*Qo�b+���d��J�#��C�a��Q#5��3�S�N�4/$�0s>W*+K��?�R�M������|/�O�4t�e&bVBn�ˢ�O��?�N�����yg�����١��P֓/�R�r`��Fe�WH�씴�W(sp�L�0s����|bu�Z���
z�_�		��T���Fr52d��a�;��T�G{�!�%��t��p�~y04q̥��f�ژ��e�2KJ�T�~��8�L�|���Z)�>�zǫӉU� ��C�0 t���qpܾ
��00Y���1Q� ��a@�20�M�4�1��^J��/������g5()J��x>�Jɣ�y���Crw�t�]���{O���+�2L�?�ke�yYI�Wߙi��$\��(�B9�.��0_��#����)lo�+�{�n����ʄK���,G Y���C��<��d�(�r�;
lJf�Y.
��UX� R�a�SY6�`��p�'��R˷��"�����Py�n 7���������]S"-B�'�RaU%d��b�Շ��F�;�b]=���.��*�1�'6�����Y�G����'[n�(ݴ]��(0V�"T�c/���/=��%pQb�%+Y���[�h鍷��a����s$@�ߍ���� ��f��"��M*ڌ<���<��$r�nO���X?$��mt� �:�0�b��;��G�s�o@�8���Q$%G�dg]�5�}��]kBl�m(�ώhBϫ�y	�Uu�1�oԼ
wQ��9�[�� �m}NT�F���:�ɠ�+�SI5ъZ�����6x�O��Z�x:9��r�4p1�)b �����
�1�"nb���� �B ��U�x��u�|?~�m��3Z���JI��x������a��Q�
���;y��;pL+����Tw�+�gbG�Ϫ&N��Н��1� �ĵ�P�I�^�y����Z��_�ԑX:XHU���n.m��p�'�I<
�&�Jm����bt��Ď�����嚌�(�7�g�ˡbڃ���L���;Ǐ;|ȵ�t���J����� ��Fx��I'�B��Z i��LcD%>����኷�^ҹ���3�ҏJU#���S,o�6��@5r_K@g�* ,�BL�a1ҵ��Yi������q��kQ �9��a-#�GUĨ|ڭ�<��)�s��#�"��!}ei�`���.��:\�-���WS~�m�h�x"s�E�{�)�]�2e��)f�z#I��N^�!�}�[���d���X���,�u��T���-����6���l3ĄRtwF��^��νM�2T+��-�z����-��ta�EQ��vDC�b��8�ca���&tu����v*1y�]F�}��J$P�4wz�����%d�I��t"����y�ID�������r�Z*���s`�ɘ����i&8�؋)���M� R,����-������e�$]`O��9u��2IZM��e�l�NiK%��95�ߤE�:�=6z����+��ڬ=ܑ��h�x7���@�W7�x̸�g�q�94k�� 1��9?$Zo�h��Ң��j��"�g�4��]���y�n�U�W|��~��*�y��)�8ppq����J��i;��P�/��eA��k�x`X��x�Ѧ�fN�椱I	�� �2~B�,8��lH�Y+�ưS�Yv �����JN>�r�/�$��I��a5��Uky�1�4��Q*�$�xZm���)���!�	�d38�|���L�z%t*�	�C���<�YUm�K�)`o�si'�}����E����`�1��X�KoM���d�_ɬnd6lzoml7xi�4.+a�;S1�L2�d���b1|VoOY�7�|.�,�_P�*�$go�S�����2�\��E�1 ښ�(��R�aV�\�x�[cVh\ĺY��L�\�HĬ��V�N���R��V��J�/�<����);�{7fS��GN|}"rc �<�_� ����3Tf@��tY�O#��|�ve3���C���0R
��A_���xb�ߖ� �=2�������'q^��&
s`��6�:���s�I?t<g�I��f+��_�fs+Q�cͺwun��ە5��1á˩���m��do�	#H�[��l���Rү�3���Cw���yﻐҗ���N �[):ޙMG鐃��s��"	C����Ƚ��Tb�����q��y�������["�Y�{�����i�
<dR����|FT(Ø9�F�� �����eeQso2T�tBe�����lK�� H0`������[���k���.&�������N���2�ڴ��~��N��m�z J�s��,2���T:�0�o[�gj��)ҿ��"m�rP=�Vc��b��%Cz֣O7~c��\Ϳo/��/*gĂ3�(W���@R�󏩩���Z�T�Y-���_��J���x���i�f'�C!n����XҲfC���z�=�¸�V��7Z��i,�7Ҷ�Sw��<��v��&�W��/wU����Z�U�Si�[�a-a`�.�����_{�-7<B�9]�
�#x�\]C2��v��؆��r�_�[�L�H��q�;Pk	U"��ۦ��Rr��bݧ��j�=��\�7P�)���qt:tM�3C�*e��R�;�&����g��׼�-)GL6/��)ޔ!=�ŪƢ����������2x�K~�Ѹ  E�Ȇ�_֧([�Mb������<�&���_�_��_$s\mj�~���?�1XB���5��S�c��;��$£����t�󑽝�Z|� IN�%���	����,Ơ�T�UR"n�l�˩��_���Bc����ֻ��� W��%9 �l���c�'�Դ�r<mA	���J���y�2�ԙ.��C���7���#v�/D���BM"�J �K�஑t'Re9��f�)1��dCi_r�@��v>�L�3��\�	���I=�~���ʻs"f+qf o'{���C�~<�]����Kg����6�_&6�[����Y�j�x�M��q���-k���oTK`���2����;I3)*�b��L��sMG�j��QB�j�6�(V�����b��ݮ�H�:P�\��{�ɐ=��e0X�G��ݒ��j��̝�u(�9���p5�O}� d$��������`
>��裄|ci��8�&���+a�H��� <��b?�H.-�2s�'Q�R\��*�*��k�>����R�����8�{���&+/��{I�u:����iVr
n����܁$��V*"�Mu1ΝƉ��{j ��mF��ܧ�*Ů���Y��2SB�ȱ�c�I��S�y{��	����A*�r�"~8ţ	���0���n�-r@A�����`�H+�?�|�XmhP�����0c�Yf�U�V�$
�[�^D���;=�.f@��}O��>�zR�F�?������Ť�����a�׻hD���^۽�;�_	�������eYYMڭ��	����׬��
��S���]��h��ELS{�ڭl0���@�@��c�9@�F������vn���=0�����ް��f� YL��An��1JCjH�RI�q��C�p��nU?C��TWZ��s��{� \�1��ү���<a��T��-�v?u���8M�Y�zO��^���(ըטPk�m!�H�q��i���n��`�{a$m��5�-�@�� �S�W��O�5]�L�/�ytSI����
��;����.W"�p�y�`������"�XP'�swv
���e�~E�(;���_�s!�]4%����Dz�a����=0���5t�����}5�i������T2��yp��Ã��+5�:��v��4>��JOM��~��1uk�Zp�v֟�-�*�[��/M��t�ٜ`� 7��]���҄����RL��M(����*yT!�P��&�]� ����"���X�߲��"�t�����My����l(h���mjU���a����l(��"�U|M}�[��j����_a�EEU�o+���v)�*�/�#�Pߐq4TІo9Ң�� ��Ʌ���l��1y`�0FL���/��k� ��H?d@}lqĔ���]Ik�OPd$M?h@��'�!�C��Q:�-��B7l�_�6�x:��>�h�0a��5M��ׯR�������\.19������uӔ����(W&��L��w�i5�ggU�+W|���cםj���͍5��ր���G׉=�ap�->������Mj��E�;��(�U|F�!��'a.B����#XΊ������Y~���3�/0i����W���R����\����8>�%����[kg��5�bvc'o��zhBZZ�U#ۿ��:�ﬧ��~���s�d�nI�� �[AB?%˥Yo��~��	��r��,����A/���}�f��#%�g���fԡr�dz��g��5mK��k�&��k�jiKb�˹�f�g���$�Mb��9����w�Mp�NF�An�B �ϮJ��5�����x�u[�c��/��@c�������ׄq�wz$��z�7�u��hg~�z�C)�p�7�*mv��N�x���'D$��C�s$�g�o��?��^n$�����ȣ��&`��q����;�%B�:#�p\݊����S�ąy��
LqЇZ�j���\
��Lҋ{�`��=3-��s��
ΰ�/��js���=��tW_AVGm��o���y}_����j%ZF��X�%Xa��)�:��Y�;xh�(�$��5fb�2ם�rx_S���R���8v��sw�i��W1J��q�s�ٻ�M��.㜟���mǜ�:㷭6���u� Sh��?�٧��A���R�C	oG��i� [�DrT�,�ou]�_�{2RO�X��d���K�JRW#9�9 ���J���ځasL�v�8ogrR�ڬۄ�N:ֶ;t19�E��U�&��-����MoQ614'Gn#z�tl�f��k�	���g��u��c.-��0i�/�"��j��D���c4�C�9�L^"K��y��z���X��iJ�-��)M��V�����+��L��^�awb��K2�e�Ek"#:?(��aj����.���=1�g%���?iCpჳ� q%�j��^j0�$�������PK����"�?a)Q@å�aj���+��35����3�vv����ϴ�TiA�ũTf��a8���0լ����q��D��t���xw�P&��N��c�>o�Xd ^��:%򁑽"�����"��e9�S�5I�K�LlH��I��(�7�L��'^9Q��a��N��_�g�
v[�����U�k%�܅����N��@˯<����Fg�Ȉ�=ۻc8^D�W�F�d'��Z�)-��X��-,�#��x�&~���@jj�ł+q5!���o!7�k*q~q�����hU8���|n/r�������[�{�^L���e�Ҍ�Ctj�������K��?p
���q�{4RϾ*#N���)�پ���Z���^��pJ��|���PB�^���]�����!7uU(_��6�Y����LBsr�@�+l���E$Ss�7�t���Sd��˝]y-Whl���?���H�!���-DԘ.X�:Úr�:"RM�e�k���a\�W֘w=��J����8�Sm#�([J�:.˘����NU�_6���)$���).�-D���g�����r�j�\w�g<?e���>()��(6�g��p*M���dc�X�St��j�Ez����$�$�"lsok�7�E�O��p�K<x�h1��=3��f����a�Q��q�0Bo3ɓ�20�E}<ʧ���\`�7�G�1z�w�����5�9�w<�zCآ��ez����&4�l� ?��Z�:����I9�n)����2C��_k9��_S\wȫ����H�'U`Y՜������~�u@���m^G�T�:EB���ӟ�?J��p2��2��w�4k)iU@3ə�WE�|Jv�=Y�+�B.o�26B���Tr�
s#0&��`2i`#��W�۵$��E���Ɠ�ƃ�x��c�%B�8r?Z�2c�C�?&�d � 0�ϟ����x#��X�kW�%��6bh�@5�����C���~:@`P?�+�e�9lU�C�|���dȄ>���<�`�b`���3�c�qd�-e�]�����XP���#��͕$G?�&Y��o��b�~���G}�zO���%���:��\���f��m�+F�i?p�Y��q��N��{��y�"m`9u��F����b׆w�+��W$`��k�Ԃ�3�7��h��!Q�@�1����h\~Y��q��W�/<�\v	� ��=���>� +�<K�� #���p�V��Lpf��l�1}U�,��Gj S���YM����x���e����d8%1�����a0��'����RI=�/�n�M��Ȧ�k���K���;�w����f�#�=���Љڷ�dڗW����6�����ǵ�!�2���.���64�-8�`?b,���T�\?�E�g=""�z�K�9���V0m����/��]�����T5B�\�7Q����_�%�*��s��K��������W����:Օ�6c˅�/����������ev��O�U˞o�Aw�k�]o�B���㌏	<)[�� i�Z$��u*�TR�I�3���?�����w1��P���p �Cb�RZʮ�T�%r{?R՞�7D��N��a��>6W]�D����a�z��o�鏉���q6������=ž�F��(��(B��!vK!-p��v��p%�Q� u��gP@�U4�>�I�G'��"Ѭ=K�n��+���i�&��i��wk�;I�R�p1��	8t̫Z�A�SbL ���f�̧���s1È�x�"��1���l ��OP�)��� z�}E4��
<�vߠ�t��S~��~�TvP_`�;�oA{!"x�WR8�ժV�ݤ ����*o����Ғ� �x ��	�=�<���d=�{	�n�y���e:s9��"t=�Hp�S��� ]��I���F͖���_G-�R����(gKiLx��6,W=c\<_3W.�`�sq����X�m��4�|	13O>#��͒��Z�U�I��f�_����h�G�d��U����дUv� �5�J�ͳϹ� 4�y��)9o�O�OWhc��|1�P!d�w����0�X�a	�a��)~�I<H���:᰻Pm-V��D�T fU��
��u^��{�}���g�טz`��rL�b<=v�,m��z0�a�:)z����
��8�8y��]�R�.L�A�/�OZ�5�[�	z�mI��v�C��x�6{�k�L��n��K�$A�n�װ��F�ҹ:�uAƱ'���x�i�,KIbϮ��~.N�
�jN�䊻��0zEc$�^,�>������0�%���Ls��~Z|9>� ;�r׿y:��������=�o��Uh=��uF3���br��_ʲ	H�m��7�	����8M���;������s�9�;�a%�j��G*s�Spg҆	4_�Ꚍ"�;�vIu�؆0�4^u��6�'H���K�K`ĨW�fU�������6 ����9[oN�A���霜����'�:)���o�h��^�I
�F����V��"�ܐ�=
g?a�Y�ڷpw��ʩ��6}���n���j��'ݯ�7ӂ[�8kM���q�F��u��
-0��[�D�������j>������1�JLP�����w�yb�۽\^m����k,�M�J�0br�6���Z���ni,��Ћ5��y
�;����ʄ[����ʴ���~����ԇ�֞22�W�⤵s��al�>��j�l����R�N�܍Q������4��bl{�Hu���&�&��%˨�,YU/0�ބ�j���tF�v��
�`�{�JXǺ>����v�*�
(ٌV�xM��oû��_s���D��݊v�����Ӂ������|���a#+�{�w�	^0�
�(��D� -�b�N�%��E�L�P���zI�`����T�G?*�n���������_L3L
�m����eK"�yQa�v�k%S����_D}������&}c�L������m&�h�����.�I{z���W���GRS�(ɭ��aP��P�`T>��jcZ�/S�Jҭl�rq�����F?�Ns0�����E?}��AAȊ��N��w�k��#l� �Cx���;��.�0������Z�7`�vב���H�`��A i˩PD{�h9���>r����$�H��Љ�Q�RĦԴl5
G��I�G{(�ppg��fi��?��Fvl�Y�ID�9��>���o'�\��NfԴ�+�ធ�+DV�pA��#r��\S�
�u��m"�,�J w�2m��0a���� �f#Rf� 	�J�F��<�S^�����Z�J+��q��!,�|ՠ⦋�\����Qi6G,I���x!�.b3�����Q�!w�
#]��>H�=q�*Bn6�zۊ�e*0x�4҄�$�`���©]��Gr���z��v��������J�d>7�	�%�bj��l��ٲ����	�E�ں�?\�ˤc�I���(z/�#����� we�B]����X�RU@"�~fVd؝����8ʔ��[�$M�E����u��Q£H�m��ŕ�[M�:%�l=u�E.����Kq�~�I1����s�&�E�!�T�`�N�T
��4p�$A��D��r�p���6� ��ed�b���gH������p~�q�v����S�kɖO�Ĩ�tp��e�W(%�m2�_����ʵ�5s��=>5,�	�G�E]J��-7�y�jA@SS�!YS�K�Td�ĺ	D�Yқ (������&�9���j_�7v���w,z�yvO5�Q�������Ƥ��T �`G.�%��3�R��-�M��;p����p��J��՝U��ц!7��g:BJž˚6�%U�|�&����U_\�i����A�D�4���&ڿ������f`~@k�a����8£+�>����g���^T�Z'�*��#U�#���?�Q|�YwO���������3�=,�ϥ �l{��$jE��m�q��^�M�'⏃�w��8�Lf���=��i�Vk�F�ezI[VO�B$��.GRׯ\ö����ۡ���m���x��eZ}B���Op/����,�oh���e������Q���Ss|��ӒU
�
Ej�M�3�l8���5]����h�]#�c��E"b$a���p@�;�n�I<�t\�������X�������$����;��i^��=
6�G�1?�t�`��^��N�: ��[cm����s�1���h<J�[_w �"�ŬãS�:� V���)\%�R Q ��2Y�S�Ԛ�4�*R	e�*�O&6���<�{��&+���p*�U�e����^����&!�ѾC����e�����V#}��	~��a9�	ұ�#jho�:�e����%���}�]���z�@U�6)����8wC�|'��9h�~l� �3������ɖH�?ӷ�ɥ���~���.�Y�*4���Y�~��ݽ�)�
�l:Y�/^ގP)��|+� lΝ�e�(I�
� >\MD�!��i�Ӥ'31˾U�ND���^��z��.!и�*���CNZjP9g�8����Jmqq�-F"�#|�.���WWt�O�^H����/>��6d"!��+@$U�R��ֳ�w3�.B��2���g����}O�{$�я�]=b,���a�iWŁ�r��x�Vˊ[�.�?��ֆ��
�'�VB /��1`'?k�4	Rw�uK�:s+D]�!zI�J|CK�D��b�FE��]���H�0 �o\�d�lw��9#h�a_�������|��B�g�~���T�������e�� FkA}���GI�����#H��Cſ<��H�_'�4}.%M謓,���? P
��BBa8�������3Ŀ�Ӱ� Ǩ�U�щ��.+%�	��.djH��iQ-����"������%��D�.vft�Ţ"5��X�!�W�^|{A���������﻽~PqӠ�w\^���؛��!�5BT{8���b$�F����^_{��ӶX؊`�Z(� !��R��W\"Q�!$;��Ζ��dX'p4Zx����7zm�ۗ'�H�~�K/-���7L��? �pm�/�6�d���b����/P)%C�N����)��&=��n|�?��ة��k-�0���fv���{,�:�@�MYނiJ#�V��n�o74$���c@w�'tsǆ0IR���$og[n\[k�+7Vx�< �G���2����8\�n����ѱǋ4zr_�u8�\Wq��f����E;&k�JJ�\3/	�\ڠ�ɞ�y�6��<Ր"1@?b��Vn��d�"�g��i�h����F���E'��[�u"���CS���y�����?��A��^ԿTi���	�������
]S@k=��dй-U$��/��=�1�N��Kx�����k����Jr�P��.L�#�W{H!@	/N�I-���F���J7�;������y��/pۭd�q�k2���	](���a�I�6y�d�ձ�B��>�(��o^=r��?�0�1�Ԡ����j$�U5Tp�&�L�k�]��ۑ�]��L��"SA�����g��!�oW>��geTz���h��t"@d�ؙ~�W�@N#���V�Z�L�'�_z& �i#��"25'�)�y8�s�y鬒V�E�d���Z���\�Te	{���@�;K-���m�%�_��Ry����^�վ㑉i,8��`i63I�Hۜ����;V��2� ��;	�Þ���0L�0연�K���cd��^��{��5ǥ�٥t����F�Q�1q(ʘ�w�1	
p��S��8� 4~f�6�	H3����G�O״;P��N�=6���%����F���ƭ�;��_����(� �f�|�u9����1��'Mw�i��ܔ�Ѣ�	�Y��J������q��s��^�Q���ݨ2-C����:�`]�4��!v��EV��)Zl|��d�b6n�=�5��Ɖ鐟r���н��Y�r.�1ɧ\��-��b�T
�,�h�Cd�^�.~�[���{_�ݢȖ�<:Ao6���"�x�k�f�8���^�IhM�l9:�����;yH%W���Ў��a�t����k�Aow�ߘ��&�S�C��v���uY�G��l`��i�Rf��{��^�F�Eq�΍.���щezp��ri(L�� ���.�u;��������l}�<��p������ĝ'qRɥ�xJƮ�:�.(�L���}*��LC��Ψ�OPkq{�e��C�Ng�ƌ�\&0=��Ӱ�oX��U��ӫIǯxO@*���,���;Y%�N�U �]�� �ˉ.�\M9/r�Q�Sz�V��w������P�Y�|����z��.��T2>����D�Ezl�ЮZ>������lBK��u���_�s��F��\��#ބ�`�������&��Kz25�ou_�T�G˾����7_��h�4J$�'�b�C�5��3��
�'�!�R?9;����f�{��%��?�D��A���H2�5[����r;��ҕk@���F]�st�Cs�;yK`h�����İ=��������Ni�$�����2���A,N5"�6[�ȴ�553�T�}��
C�Y���%LӮ���4��Ӝ�[{;�rȵ�N�?t��h���V��/N�.��i�垇6�rjD����Vc�]��#\v;W��З��7�!,ʃ�9:�-���4�����+�j����H�4�e�v��B�C+3n�adA-i;�;k��6(��D➘Knk��0���qF��"K�rA��b\v9�����!�%M�����65[1��jpk�)&�ȃ�\>l�0�d|��͎GWE�p|>Yh��봶�P�DG�DA9�.�@�h�����&I�M���7���W}��<կ��H�Qc���!�õ���s{\��{�<��J�5(�E������"�5Fw5>��7bx���`�vz�-�%�����=m�O�7�Jo]ݜ<��H͹�+�aɶ���?�Ȑ��� ��k�B�lE�g�N�gSΟ@}ѳT�k(��4��O��K��_�Ȕ�<�~��'��J�H~���@��wl�n�2�<~%�J�$iy����|V绱���~���p�<��c��fN��fs!8��IBn�ޒ'LR���z����F����Q�4b*$�/;�|x�j��-J3ycĒ>����cOd��6���F�Tn>	/���-����Z��#!�)Q* t1_O�}�h����Oi�4J�F�.2��uo�.��*�H�
#q@��WU d�|%0�i'�[ !^�x�z5IIh�ZSy����*��>6C'�I�2ރ�J`YG	����lum�b��F��}�禇���k�`�������	25���T��'2���=�J����~;���.rI�jGOQM��7� ��<�f{[��(���S��`h�AfsD����-n�N���irpO��s�˙6|5@��ܶ8��/����L�F����4�X��ܺ��j'���v�kX�(�L��؄k��?z�s�L�J�#��Y�rƎ|�N�JI�9��+V��e���_«�W��:��6��U�V�[�j�����MVC��v���l��1�BK҉���OLZ ��w��9�Hޟ��U�,�B{��O��+5���X���B��(d���t/����T��設d�=#�T�ayV�]'��/w$#��x��ɡ�$��x�i9�[o��e���ǫ�P�e���I���U�����^�����1�1�O��1��/������챼�h	�}�@5���nґ/��Z��v�`,X}�+� k(z{�Ѯ�qK��l;�.�G
MQ����VZW�k#�x�}�n3E�?(�3�d�/8�o�h��	�p9V�ĸF��/�9�Kj����Cl)��@��e���T6j��2�j5Ӳ�1�=���b]��}|=V��x��U�'��_�q��f�vⴭ���5�2�E��+;XX x���=D8�����%�l:�GI����Z����Of���↟�b�H� �!�ڊx������π�>�j���c.�I�V��Z�t��

1#��Vo-:~^�~5;/>�>�y����u�8QP4;:�^7���r�!���2�O0�-��`Kx��	�9B�W�֒�������7y���sXF��:��F���{2oP���"*;�ߋk�E�P�{M}`Χy����퇘n�5�Ēf
'�;1�
|�x] �_�X�'���YzHC�:߮��VtcP�\x(Y�g����$���h�ədkH�L�C�5���vh~���R���*~�b�T�3������|�C���pTD	,�����b�b�'t���Yv&G�Xe7�D�u�Ӏ&h?���t�ġ�z)��i2��Ӄ��;�P�@���F��˰�n�;���}|�a�2x v�����Y���4NZ�����	\4R/:���i��e����a�1��1�f]{f@z��'����c$��^�	�MDoC��"��-?:�'�[�vsqwӋ�:�+gV�#�[E)��V)3C=�O���,���U0|��s^�@��#9�A�H��WY�L�5��"���On���a>���rUC��t�(f;����nJ��gۮ��(T��9�;�t��e^�:3
�?�:��0���'�Kg�,�,*�����
���dGmj���ck�JM�`��I��Уԭ�b�x;�R�Y�SO�(.$��8���b�{�+���V�B\�mMFp�[mI�JI����;y{�T�ȼ|~w�͓_n��޲G�'�-\/�v[����G��1����"��*�~R߿s5�1�a3h��Y�\�DЂ��A�`Ш��V")�S�k~��?DH^]҇���2���۶���^#��F�c��QT�A�=��?����(r!���ֿY)�A����i����JS*n�{]T��rF��� �hM[��?y�vM�u�]����HN�J�De-������,�j��%DY� I��z��l�s����b�dR#�\�N*�����'����,��;��A��gƋ�T��y[)$�/r�E�G~UĒ�o<�B�jr�b������V�����;��I
Q���v.�8�y�Q�"Z�Uy�zޭꨝ׼@d �	ʆZ�����wޖns+hj_h\�D4��3��L�"�����m�ݹ�W]R���j�7�ۗ.�~s[,y��C�n[���J���������~��X��5��&:,���y�ˋ�<���G��\
�T���r���(���~�fTiE W.˅��7��>����B&�B/�P������=� |���a�gm߭��gB�*��!��nv��uk����A�؄�K"J�X>��Z!��Sl3U�ܕ8*�C���\ʉ��F���EEm�_�����49ߒ��v�B2X���E���+`�C�f�ߓP��Ԅ���� r{����
j%T�רZ�n�i�O�;Sɼ�����*�4Pp݌)N�i�����s�m�LA�<��$๹�v��A��[����i��UA&�\�B��{&I,r�"^��?a~�D�b
�v,)�V~i�
^t�W�<|e
���R�g}^Z��6�X�}�OdͰ�b+꡼���<A(��Y�;ڮ���t�'�?��Āy�8x��M����N8`��y�������fj>v-C��H�|�.�`?�b��M��[Nu(I�Z��{=���4ݩ��'i�Xڗ6˄[K�:`�Rد�D{6��e�ya� ~�[��+�ݲ
��-��J������
,��|�*�I�UN/dN~��u��Sh�I��-z;���p���	�[�*̛Td�Gи)xK17�G��}��(u���TH�=pxLփ4�;��ڳ�9M,��<m�_�AT+�1�q8a�9��W�-�0�X*�Y���v���{oK�=8*k�"���+/�zڽf3L���u�Ck��O��[-x).9�*gm�u�Hv!D��v�b�~:�
cP����o����#e���eԷ�0'�%�1p����~�$���@Ga�rf�7�|3��$���m�<m	-'J�ƻ�È�p��z!������3��93���Qf�[�������q\l�h�eW?�I����e�(h�zEۂ5d�_O1wȌ�N+2E�V��8O�������q�:��z/�'B����d���Q�E����?��@W�s��L{����uLg�j6?�a��)�.���[ۻY�&a!s1�]7[�<���^��>5��;4;���ZE�����'>(gW�lvj��v�������n_��=���r��t�V��W����Q!��Nz	0׵X�o~��3P��7 &T(p�I��ٞ���3g��sS�3�41���J����C�e9��A�i�m�y D���qV�Y��C�V4VʁO���l�m�,J���Ck��R���ʧ�Ī�~)���𽭂��r�yT��? ��br���!Q�RD�L�)Ze8AS.�`���#��M��\�щ���5)�3�S��#��p���w,Ho���Kz�egB�Ə�H|��獥�^�r?)���P�;�ZK"�a�V�MKn	�Xr�&�N��4,�Y�f�9���$�P�%1:�\w�U��'$:����<�N��|����h6^&ˈl��
/=�W-b@��1>��H>V!��F�gۧb!Ԅ�2��"�J�y��ec����O8v+����*��[L�u����uB�L�m�΁'�&.>K#ȼq�!��'K:��&�@ӌɤ�pu�e^�9����<���O�����qV*d��.��`l�>R�`��o^5��]�h5����À�wTWJ�߰79���3a�X�Q!c����C�/O��(O�J�[�� ��M�
��!�m
�m�x%H����q�1���=�<eÃr��Ʋ�mO�Gˆ�_T�!�b�h�)���2k^�Q�Z����L�m90��{���Q���Q�}_H�vQ�G�O���{0������g5`���>�$��;C+O���^�mU�������ޟ`�,�1�=Ʈ�.�MD��Ⱥ�<I��
�����XZ��#lf�֌c�� �z�5��*�Pe�jT�ddZ!<5��b֌V}jG��-�.��ݫ�_Q���N�rzcSL ��T(�
+Q�^]��<�v �T͞���1�L �n��X���}&1,&����K:�#
/v�P��H����X{0%F�V�������֏[v0�H@q�x�ңi	>@�.v�S��9��`~(X�?��D�Yv���g@x���{��1��-g�]A��OͲ�LW ���5sۚ�8۰���=���;��,��/r�Nn"ܒ��t�j�~6��&�	�j��2������ .%��b�ȵ�����@����f@<���W�S��Qھ���x$����eX,�0OV6=��+��7�Sq�Y��շQ���_ý_#����6aߊ����1%ܿ�R��W�:�w�j��&i[mҠ/��UG�,v�`���1�5:���U�����|����*5�_zQ�f�Ɂ�p۞�,J^�S3fyɸ���3;X_��J}>�L���[z�:?3��鏹���V���y7ޭ�u��`�p���*���B$WnK\�8:�p<Ы�1o5�#�OK��c����e�[�fũ���m��?�g�?nk��� MC����؁U*�/��.��n�������\.��4���F� ΰ��v��˕b�W{�둦����.t��$0n��6��y*�C�奫�h�`��EE�"ޑ�Bπ��=���x�HZ�fu���>q�i�8�"����և3���Y���N����k�׊�<�����6�ĔޏA��J�ꔳ�w�Z�&�5}A�J��Y]�J��~C+�J��(%�73ؔxMU|QZ���m.�c�c����ݐ��I�����Q[�V�	1�[�3YgQzpQ�:s17�& QӅ;C�#�$�����w[,��B{�K��d��B]L̛J>�3��,j����L��`60� �w)*?��.�:\��T������.n��F*������*Нi��w�	���8z��N��)�=Ĩ���~���ݐ_q�����>������.m��ɥ�0u?�iݡ��U	���F������$#v�b�`�DÑ��`�O��Mu�@t9/6��=76[��о�����\��Ϭ�ȶWn3���>.�K5,�&��S �dהV}�ϲ�L��h�s&��S��U��a���w�n��r@�"Mv�f���@�t
�bR*�<Q���&�.:]���K}P�P�Qܩ.]Ү�9��d�D���N�B�F?;�� ��{���g7���d�.ْ1�Ak�ͩ�! m?r��8�1 ��Hz�#v�b�/]�*r��bE�@���:ȊJ��_�\��[$�1���q����Ҩc�<�?��
2K������%ڇ1�����"k�X�:�H�B�@K������_"5S �:%��z�˷6�g߯%T�1�6Y��Q4��1q����m�F@�ϋ�������!"���T�^�YvLH°7(cȣ�+»SXH<f�������-��
A���,5�楑��8Q��]ظ���ѳ�NZ��i�=�����M����P8R�N����qs7j�c���=�����UTX8K#�DS5E���ڧ=�k�V߃q�+�g��??ńTS��YD���J��#؉����٢���;�Jp�d7d&�����9��n���̍����L��Yt
Y-�:��b@:?�1�ޝ����Ά�݇X⹉���M�BF��p���%�������/e�Ћ�TW�	�TQ�^�P�ˤfA���~4��~4�� &��� 7,��Ze؈�`����$J���ռN�O�zU��S0[�_5�ߢ��Թ����C���2����,k�2w��>�]�ol��#@�U�f��]5i|���j>7�FiyIe(zhmNhEQߘ�$��x�
T@T����0A3j�<�},�0�c>.�W��:$} ���z��n<D�7�8}x�q�^e��2��W�����17ơ~�뙑���%��6�8��?��)�{}&DG�Vg���I ��4�YwA�A,�ϒSX�I��j*V:_uPȄ _�#�n�$�fp�\�N����!��zf)�zW�L�k7����"��&1�NSo�Z�軖[��Ĥ�%��Vl��|nk]F���~4V~�ގ�͒�?����p�̃F�}IX8�z�4�}����\�3��Q��	�kbP��/۴�ʌ&���HB�ꦵ4��=̧]u�M���`�%�4ߎ�A��s����V�8����F�/���w��YLNFԚ���o%Q`�+�|����6����8f���Ӓ�U�Ix���G�à��۔�S`�UՀ U�H�L�^@@?e����_�F�QE&bj����/׎*�Zi=��m�Hz�-��j�!ia64�/VM[]c�6������%1���gMRE�'�K�XӪ�,�Q�sr?k�an����qX!�s�>��u2ܫE9�1V��Q[W�is���g�Yj��l�v���/.���x@���<��C�0�n՜W�����F��C��$I	E�%�n�rrm���z��d l�Z`"OƪԺ��M,.�Q�Q?o��eSFn�ᏃBW�6����:3ĸ�(��+b�=s��Ӧr���0��C��ڢ��N�Ew׉{�.L�׷ɸ�o���q���[@����8��8i��6c���+�0�X��Y]30����),4���<������@$���'[�����>q@���.�j��*�� ,@�4"B�dG�ն)�No[�-xb��h����U�{Hb)�x�a�"�[��rR$(��H`2�^�ׁ9����M�����c}�Q��Cn-�l�VK,&9��L1ڕ�"��I�Y��0�y���V!�յg�ѯ�I./��_\��/��Ŵ�3��^���z��\T-���U��[���_���N�Pڏ�Ez�p�bݕEGyt��	�	���o��Q}���X'b0�?���A��Q�����%�-�مno�c�X,���hb��$83�D*���D��Z��:�~�P�J��kD-O˝
���'pD����$!��@L Vm:��$��7���NJ�S1.�;'`yԱp�1YI������V'tw���+q����������~���mN�/�q�.o���#xG,��' ��r����|P@��q�k���2��q�%I gN+��	K���GE7�g�������Cu���.M�'K���R�j�Ǚ؆Jׄ�l4Q%
��Ը�b�UUK��4j)d��n�-���(�>���=Px8V���O%����2��A�BV�N�jiʁc��}Y&�<+�䌖������TMU�˔�(>�΃N쫚סwL����$�x��:F+������,>U�t [GLSFx��D��S�m~���oQ��}^��E/�b
>s��y��WȾ��#�cz5���E�,�c�z�(�w�����)��z��������3A=�᳃i���_Km��/���g^`zqa�-k���:����]O<�������pgܙ�ù�\�R��BG�q?[5UGc[�ݬ�}�B��R�_�_Հ� /�`�����6&�����.�k;��b��̒5�N���HȪ�l����E��%ɔ�A��VY���ٽ�dj��RJ~�-�S�j+�lQ牏���b;��Ӿ7��Z-|☲kj��cs�Zx�i�:����/�=���5��ʡ��e�DwG*jO��M�[ξ�b�Q
��=p=��f���\ ��>�R�Tz�G�\g��R�5��ʖ��xȖn&���Y�^J��P�L��fy��7$�!�c�U����8y�}�E@a���_�!t�>���@�����
���j~���.�]�zS�H��:�s�S�)c�P��*f�Ƒ^б�#9��n
����m�/���:����4��Z�����7Ih�ϵ� c_OxփU�))+���!��L�l�,�9���R]m���6�EE�xS�jm��N��@�Rvb�+�M��,�.5�ď�J�G?��9��K�q~fl��t��#��74qC=�o|v���7L��8v���D���N�K�O# �cRQ>�ͺCĀ�l��0V�"�O���h����c_:gk���MB.��k��ږ�P�W�'�5�ߝ8f��Quy��S��Q�O"Zr�e�U;GW���A�3�r�cp\2��Ou���'����~��׷u���m=��<IW:TO|'���P��>J^�: ��<̈́�p��hs���Fu�}ݕ��Ax���V�q��P�Ȳ���b| �%S�U���h��x0�'c�� z��1Wp�/j`���iEw6+�!~��٧¹i��6�J�����Qt�/�&�bH(�JO��1�Lѧ�r���;�ѿ��ga+Y�� �a���$���D�F�r��"w͖�ǖ.m�=��yn���Q��	u���f����!���j.t��&�M��� x�Un�4Ke<O� �F����U}����+a��� Dp�(��d����N�}gd�c7�c�K��fUiF��
1�W�C1ks^�����enfz5sx�;� �̞M$%T���s@>���G9�FonP�8ɍ���ja���ְ^Is���@�3`'uR@�
{��9��ތ0�i�����FN��+ق�V�w���Z-��v��.��N>�ͻدk�y�@ �o��]F3%~�,��4��ِg$�'���Q�5�J�>F���S۴�������7V�B�l5HH�*�qd��@���تAaC㝈���s�(?t�7\"8�ڛ�ۤq�-�V�\��굄�K6Hk�5��}Ķ��1�ײ��}���^)V��@z��F�fɣ���N:18�("����ډ=3C�W���Pp����l=eWj�y���-j.�7��*�����pg�z]��)ׄ�A�D SPw�sz�x��mt'B�E|�i����94���in��:1����^��Qbr9G^����:���J���?�Q�l��Ɉ0��kf�[���?m�i�x+��O����r@��x��"���zG}�n�6δ�1;��Cz�Nq�S���x����SN�jXù��m�X�.�A\̚�*����/*�W�0��!��(�}��Z�ǀ;�ώ�;4�Ţ N炜<�����G��*ݐ/��#��D߰ ��_�7͚��Q��@�nݑsx�������¼?�\��)/��@v��Q.��Їw�.�I��&A������%-��)L�T�t}[�:p)�(�D���l����J��Y�%�L��I����k*I( �6�Q�٫���I �����b]Yb<p��%���[���R䚪�c��&&�c'�L��-1fOPb0R�}��>�a{d{�����Y��'�vD-hE�خJ"`�v��ۉ���bDT��P+=c���R��Y�����b�j���)��`R�;6�^��j�� ��;�����K�-����q7-QiL��K�I0C�,�Ց�	��;���D�(��*�8t���rR����C�
�����5�'Fb�n�r'w�ɛ�r���}Dv7GԿ���/
�Z3e���}?J�`tU�� �i&4�\1��k��]_��۰�|�ֿ��paT��O��y<�Pe��&���C�餻�݃�8�p}�~��$��*��w8��O����B-��ǣ�_��1#��0�Y9}��Ʃ�=�ސ��F��Z�@]�����W��~���"�Kg�Eza�f������Gu�/��M(&V��F�c	pK�F�\�u�%Y���	Wo2Lڞ�>�D@(+���{�\̲L�I�D-p?�m�Ac"���Ѱ'��7j���s	��@���+�8�X�����vA W#W
������ר�����Ɯ��I�k���(��,�_�/IPŹ�@�\c�8���:����T�8q��H�ˠ*�����j�0���ٝO���Þ�Q�#&��jcڮ�s�&�j�D�P�( ry`��ai1QO��}�)����kr�B6�O���6�=-W�q<o�[֘ҕ��U���,f��z��m;O�+L����RJTAR�3
�ը����ܞFe��/��V����	o���*�^N��v�4�I�E�2N��`P��N��Ɲ3CŊ3��ʙw1�M�~�h
�ݒ>I��3�C<��-�y���%����[�z���M#�����K����8N2m�~�E���R��2����J���i��3&4p��1�U)���ث���R`����!W�$��d(��u/xu�:Pѡ��Z͇i� HY	���Z���T�	b^�皫C�ľ.��j�܏�*�����W�����C!&CxOC]���j��}@���McmM�����Tti�)W��>��ěG�zl�<RN�]]N#�$� �u�M���Q�<�=��Z�f67��:�E[*��C_5�^�@��Me65Tǩ�m*L�\�Kz�7xN�?C���x~�I�Uo�;�K%Cp;�z��������a3��	�+[$t�����Z�x�M�Q_QXh�G�c�\��ë� T�VpH��rofgQ�O!#��=v!N�?��_cj���;�v{ ����6�
$����F����~����<�hUg�o)r���נ<E�TY痷��Zf9���	f�ƁM��1�GR�M$�����yڳ��UL�ȓ�a	���pt?q�~{�ģ5XH_1��L� �`��K�V�P�MJ���~��j�а/��B�H�y	wq}eD�0`aF�Y���m<�Q,����ه���w��Ε/:��y�(��%3b�u#���q�\���n]�����n��l�\��W�TZe���$h�D�8!ᜯ���&�a���L)Lŗ-�k�'��>�+<�����,��PjWk�<b�@Ub]���O�|�ŲQZ1.�;�������T���p��}�$>���4�0���K����e6���`�7�}K9���b��8Һ�@��a���*��i� ?�m*�W���r�$fx���R�9���0���c��GW�v�sM��{�u���Mձ�d��)�U�����gng���,��!�pK?��HW���4�r���#��m�]/x�h`����P��=� ��L�X1���>G=FE�Wh�ԍ�2W>�K�/�R�\H�����~G�.�8{��Ӹ����<��p��q&5��iQM�}�ҺCt�`�}qPx�7]��ߗ�B�f�3	���S��}`ۣ�X�_A��KkD��=QV�����|�p��k�f.���j��8[9&�Z��h��*[Ԉ���U�����s`;4��/(��|=@y;41�Q$7� p ���A���"�╬V��p��̠��tG�V!x�)[���y~X�\���,u Ő�O4� >^�L�f\)�����LA$ J�\���y����~nH�WŘ�.iђ��mǕv�f,l�=zdX,wŤ��ROCB�$8�>�+�+'�x�O��%�".���-؀l{fqF-F����bD88�4Y�Ao4g�W3�	j�xV�h�����)�(�������|� �Su�:�){nT����s6��<~��?��/���W��^�u%��Q�}H��y����]�]�e�bT9W��~�f�$�D*�AY,r9��ê*�"g��f1<�H�0� �w���'Cp(�j7�*����}����*��x0G|�@�>��LXc�����-_�
����V[�Q����&��
�;Wb�ONb�>;y�5iӻQ����~HS�OKWt*�#���˩m��x�Q�U�l��5��]��&�Rp^��b+�:"�b�g?���I|ݗ�Pemh�z�#q
�͙0�qyNO�@3��������t|�U��^|���0��9m�$�X��n������CW���'v��:�u7�EEF����'ٗ���=+L�����N�i�h.٘���h�A�m,�	[�F���FBL2�I�lp�������	�v`�5Cfr�e�K4�������vN+�{I� �B=1(�f��=	�+�Ɍ%f�*E$Ь����c����������
���$�9Q�d��H�y��}�QDi�A���՜����k�=�Y��
��ٚ'�D��8�v�Փ��de� �'���e)��ۓ��(�oØ~�I����ӈ��{\��7���Ck��y�\�^���������A����`y߲���>?5Nz~_�>���m7ޅ�N��oI�~&. $Ѥ����(�DȰ�lZ�K����%���5t�u�h_l�Y�T��;[�?$d]1�c���,�ax$b80�[��ֳ^�������ēQ��in��U�H_������=�	��Ҷ��t�R���dv��'������0�h#�u�t�IX!���57cj�G���(r��ĝ!�_s��������k�f�Sf��E��;�� ��>��0��F�]]��1W�-?�c���/��:�o�x3�G���F>�e�<o���a�3��A����7+��%C72�>�H�����p'1�vښ)�uM9XzgQ�*��=y�\b�$���	��qRs�G����D�d�=$S�5ē�}�B��x&<��ia8�zBU���(�ƒXYʩ������t�%�L( ���]%��A��N�vS�&||�@d8�K�, �$��Z�w�l��[c����u�L��:Y��_�J��܏�R!�|qgk��T��W�MbQe���)�t���z0��s��Q	K�y6S�W¾��~_eB�g�=X��Bl�X~����O�fޓn�1�Jk(Ԛ\�\g�g/P7n�̘1�y�������l: �3M������Գ��?�n�q��V~���ob}M���6AP"�"a�$��t�*F��i�U��I1��s�"k�r�d��7b�l�T���.�'Re-���>1��>�%��=���h�a|�DՇ5�pLf��W]���x��Sj9��}���4m��e�J,��Y��{����E���z��zsֽ�F�.Mp��}H`�ܘ.�R��+3.<d\���&ލk@��_k���-��)�r莶�2�J��bA,'�8}!���1��'ҏ��˨pQ���T����&��݇c�L��X8]N��$�,/��13~|q�^�`E|��9-9�T^=��2�\R���g�ķ]�!�ͽ��Vt����o���Q�ql,3���4P=�:n��i
��r[$�ok��J�p�ht���3:�H��uu�@���v:� �,g�J��^�9���8�'��?����T�'��׻B���lґ���� �ߜ���h�Q�f�Ѣ��B��asQT����~�H��Q�q��2���Ȯ�Xp��p9����]Q��'FL}��{��@��"6ޒ��V�㜉�	�I�oP���j@Vk8a�7�~#�Ny���rl�`� �2\2��D��n��(Q�q(I�aҳ�e��cU�X�rڜ�	��F���Re�}B��V2��:Kq0x�p���y��jaڈ�-1
�5v>��ȚߢI�?LTS�Wݜ��@�9?���A�ZR��G�bi4V�� #�ʿ]R��{��@$U�e[�}���dXOx �Y�+.#6�d��^O�يAVx��s�&,.[p1w�`��k�:ZS��,Ln��|{᢯�Qȷ訮�؆.��@m�_�ŵ,B���c�����E���=9d�U���3kH;�������k�u,�*�ц�\N1�ڗ�|�[:jP�PԵ�N��>�%�������ד퍁(ɏ�4�=�1˻qB�B+��I}����k'�������Gzza���9������y��'W�Hܟ�.v�v*TT�a�5i���X|h��%�	��x�:�9�)�le9�e����WT%),���H��"�<+�P��>������ǎ�*����0�6��3�
��{6�Vk����]h��ޝ�=УW�~ǵ���y�j )�{���ꙡ�
��+������4�Dq�;f6�*:�q-�h�k�D\�X5�1���T.u����������W!�$��P�h�6{�LI;�v����8�m6��`��U�>���L+&N�����8sL�\V"�uG�� �+��!���c��V��]��=����]P��_���#�tk�&����?Q���������p4��0 On��j�������:�����N޹�c�!N-P�_x�C#�Z8����S�h&.
.�!�}��I����(!�xcܗsȴ���#*�R�BA-����̠�m�v:A��M���ѕ�C6<�JFT�⑄�p�]�t�]���D��#���?�B nd�����5��?��>q�����(�K�M��������a/�I')SO�_�Ș��
xO�E�����KI�7�F�Y��ش��!,&CQ��h��@hX/Ѭ��v:3q��ۼ�a>�[��]��[���:�':p��E�"p7Ʌa|?h�G�n�h�6#��nR�e�I�|D���P�*�$`D�	3�&Q�d)fl`ː��W~����U�״�~<0𤞲<��h���N�`:C��lbZ"��(��K���Kz�:G~�P��_�HM*�L�3�ZE���5'��<�k���t�}�,:��ݰ*��;��M�����\��*\�v����[�}����:#���ʹLY�����p~��"f����Eh�c��Ącj�dֳ_ۭ�C�����UƦ"���A�=�\^s�>Y~&����a;,R��3ms?'?�2�V����7��MTD�N��ɼ�Δ���Z�G34vM����)�ե��t�ѸM�|�{�B�̞�&�=����}�- .�]��K���~HIX�%6:M<��BH��H�vJ����ܳ~��F��5q���ߡu ��
GVx�L��������B���<���מ}�>�����`(txi�J ��)쩃���$D���P���\� ��l��!��&R)qא���gv� H-b!v!�1�(����+���B|R�E1�1�{�9e�M�������1QӁKj�"b-	$�:J�{�Ο�#�h�lCZ�/^��s,�}٤إ%l����h�'��"}Lw�t�|!qٜ��0��#a*� �Ss��  #V�����f$B���������w�Kh�rMp�K��ϖ��QV��9���̿����F2�i���mB)��'���P�h3��`$o%��`:�3F�F{�S��/|�A��NQ([����74�Y!�� �F"f+.f�R����z�w�du</mH�G�W.��AWe�£�=��:�����-�i�n����f�I�uv��a\6!u�o���1��V�$�1DLPȧ�������8��̷� M�e��͠��c��w����:5���LSt��g��� ��&o���۲��:��,����!�Yf�C^�p���i$����ŉ?�]�>�5�},j�rb]mfH�j�5����m�#��elM�M�aC[���q���}�(���~X"�/ � �&C���n���lY1�E�D�����]��!�;`�a:�f��]-�/�;�"*O6,�d�Ͼ�X��zt�@�M�Hh��ׅ�$�҄�F�PԤ�{���7��
���55���̂�>$n N�h���M�'�3k�'1���BR?�w� �k�f|^�/N�RascxzkP�� ���'.e� 
}�41��-����ի�v�_��W]$XS��7�Y�l6s���wt��8nu�5�7�d����)<J��ee���~Z�|�K�W��$>¿�ұ���Պ33��ؙB<�&��#��b@�*�� G}�/�,����*ʰu��o�4��L����;��YM4�l� N�D*������0����N*y�?Ȇ
�m�j��:��L9J�5�˺w��Y�p��%����COu��C:tS�|=�n�=�.͕V�c����ܙ:Fi�3�9� 1lAU���������I�Lx�a�(���P+���6|K���
��'~25$-GIh9��G�U�4^D���/Q�������z��fj��~��D�q��@1�{N>v�4�:��t�\�B6>c�*�5P�$v�Ũ�*Ef����",(Hu��י��'�f��t�̌�t�szw��1�v�3��4��_�i2�=V (B�d|�
st0(`	�����"9]0�/�s
�S�dV���K-C�c{�u	U�s�بAn@�n��.V�q�'«���Ă�0'�B��VR���u[F�R�o������'!f�)�\�e�J��dϩ�����B��)n0bx��@,f��p��QTq��o}��ˏS,�V�*k�ab�s���<�,\��H��%�#����< F1v����r";e�˙�LI�V�	�O�>�-�X�z�~;=V��UN��A\N
�:�,Cӊ>��B���J(�2T@l��	�qi2tJ!�6�%oʔɯ�w>�Vjǡ��� g�vP�/�wHL�J)�X�ƻJ�����Ir�&*(�Ë�!�x�g�����oc�~����� 9�x9J̭��W�PY�He���c����Cǟ�H�*3`s����_m�6���d��տ�^�ۣ�(�T�|d�\XeHT�P$�XHa�J�m��'L���#+�0<�]��X(�%�ƥ!Ϻ��:�J���I)�a�Ӄ���Qҁ�2?�\J�m2�	a�hY�G�@qXj٭�8w�)��G?�d!Q�F�c�N��J{�}���Wͥ��yx��D�܇��S����}�D�������\�gc�`z*�`�+��>-���-�$�%v�	��0�mV�ާ�1�c@��T�� d"Y>���BI��l�l(.{$<��*\t;��$ac������d���es	�ɺ�U���6�6 �N�3f�����NA�b7���]ᙀ�#�>I�p+�p��h;HL�t2�D��M��8#�WO�M��&Gv���t�aHwd��� ���`I�a��
3�L[��)�w�ۜ���G�	��s�2�A����w����<�K����a���ΐ1�ڈ�!uFje�BƤ�!W�QJ��P�vGZ	r�@�ꖠ�CQ���%����&���%��۩�y�F��c�uMC4i��!��[�ݚ�z�臙��
�zf��F�A,�(�v�)�^h���Wҳ�L��E`$��Z2Ԇ`P�"yv�SK��U�A�|�f�}(�H)���-g&1��]��,�#����
�S%�A8鏰��.��1��C�;Ki�j8=��u�}���;����˛�G�J,��#eۆ��_�9y�nz|���V8����X���0�}�8��'q��V~�g���in���\�9���r�=*���7�;$��<~����l�`�Ym�2M��t�7�:�c*O�: ��c' ?����[�/M� BVms��F�o@�,T^U���6&�@?���|�T�밙�>��N���k�g#i�&����Ul�9.�xt���r/�{U��#�KF�9T@~u��K�ǩ�ZȞ��3�oA�����J?�rw� @�(�J�u���z٥s���L8�
��<���s��|2�m�J���)KQ@���<s|�Z�d6[�?b���2�o�ק��3����Y�������&wd��^���"���n��� ��y��1t����i٘=���R��tmOy��������՟6*!C���a�!!��k	|s���L�zX߲�Y���L;��C���{_J�:l���������fKO��Af-dx�"�dEo�D�:T��ŋ�{]��vgx1d��Gܙ{�����K�QL^��\O�n,�����0��M"�N�� �%{F��~r�@^o�;���Ը��2�mZh 0fo��W�%���"��A|V���fN�:��|9�+�>3Θ �M ��T/���q��%�uW���������F70�	_�f%
����z"-e<?N6'q�>�ڿ\��v�f�;�[%��hh�t��"fvs�7������ߜ<�gW\�ȫ�o�F\��:�]u�c�t �HԚn=�%����G���Ⱥt�ҳQlRl��:$@���-��A�c+���f5��u�F��_���ڻ�2�c#���#���9�:u�>�i�/��8�:[�6os���U�호�p�Pj�V^��}�s���:�wK�M1O&�u��.k�w���8�˼��FB�KN��%���xz�~x{�q�_���M>G���/�H�<��Q�Fg���>�~l��=�����5���ߍ��!1A��U�b�'z.γ�F�����m&
_"\��A��[�	R���[�'���-czðN�PR6�Oz���B���2Sۭgv)>�FX�y�:f��&�&�2�)J��}_�n���Y�$�8]�/jE�ų�֫�S:^��Y�L&��u��A1�^�@�`�տt�8o	�]v}N!?�:�|��U؇i�PO+�eY�{Q��	�Ko���M��!ѿ�36��+�:�O�ɭ���y�|�z.G�E?�g4:4cۮ��#䎕�9�M�#`�"4.Q�
�������d]�!���F��ǿ0
Z�u�A���A�F"�m�C���۬��<h���0�J�X�nQ���@d���:�_i
��G\I0���g1�_�~%�Tx(B���sڌb�N�+%����\�)+�3���桊��V
�O����c��Qk���{/�'��0�,fƇ"�JC ����j�>d�o٧u��T�3U� `�@ƯYض0ӿ�ɠuw$Z;�u���f�9E&Vߥj�`~�zm};�� \*s��=[V���h�	兎�C�^D�Cz�-�6�z��arTQ8�%�䵀[�)�n��4_���A0�`SXb��{����Q��e���Ql73�r��>��I<��ޞ ��Z��d��8\� ������S�`��9�9l���)F��Ua|���+a?��Y!=�Kl�8{^�[��^�R#�1�����(�GhQ���ccg2
o�(.w�`uv�;���w�h��T�%�hE+�f��*T-���&��k�*��6����)���<��#%�E�7� ������3ә��2t*@��袣Y�Ǣ��'��Q��Ao���,�b�>�5�hw.*b��&F��З�Et�7�)\��{$�?��՟���F�N�Rp�.μ��S�v?x1r��@T�v���2D/�r=9���E��}�2��.'��˾SI�"C1��Ȫ����{S��<N�k]8����r��J4W������˴��o�ի�pջO�%Xj��߮��g�x_�*S��?�B�\�S7	��oi��	Ar	2��Q�*�E� �H)*�{�	-��h�(~CCB������5��}	�щA��	TG�Ej�����J{��0.�&�Ng�7Ii��^0�A��x���)����[�F��Qv����({6��L^�.��3�=/�\^��7�Z�o���U�lh�_�Q"���������%�b���Q��B�X��l��v�?���#��q�Ҕ�1�"E�u�)�"��yw_��BW�d�
���������nH��^�#��4�C�F 0I,Kom
�>�I�,�:a��|�reD�+A�mf������zn*�&	����&~���8�v�ZT�~	[粿u۠��yBrZ���!e�I���?�"q˩ģ���#�D���-QҰ:hq�T���Y�9�P�z�!�:_,�)+���1v��72�}��z���X�B�ٱ��}(�m��6]=`Ǚ~��S�Qp�Jt[P��ll�w�I�iRv"�A9�9EϷ"�V����HxTQ#J��r,�..#��0�����%�F���]���9�|�N
k:+e�QB�Z����3�x^_%K5�Ra��v�NQ����(�u+Ɖ��K�W\|�*��rkg���O��զڧĩ�$f���b9r��,h@����#X���Iy��+Λ�����e��a,��o�DP��vLI�Hw��g�d
��@J'M�Vr���ί���Aq��N�ߐJE�Lן≠￨Bs�fo�����������_�����T���}k?(�{�8��~_���=�.V�Ŷv��]�/�D�g�X��5�%N׀R��N�>l]��Ŷ�l��� �c{f?�����P�5�d�m]T�HCh�E��$��௰Ii����Hj-;���VB��;���B��ݡ�TJm�]�:�f���|+&}<����R&����92P��I�����$D8K�4G d��3<� (��j��B/�ꭠ�`��QN�瞍�$�F�m�t���a@��|W�9�:岊Q���H�^��*(�@�3�����((�3�M������m:u.�iW:.ǘ����=<��+�d%3r�����U?�>wǫ�+<&P*0,���Ac��.���z���i��w�]�[u�M"�g���8e�nPx����Zd5w7��v�Q@����=.t�+]<x��$���%�s�*�ӳ7�.ȷ�c��V�,Y^*S�"���ج6�t�w�@��������,��(��{������Sm"�ڋp��^+�{"�����zOe@�r����累E���(Ɯ}�����뤨w.��� �X��b��=7_��Ly���G�o
7iп��r�-V" O�u�ȣ�oLA�ߋ	3BΦ�n@Wy��ҍ��5�s� |�^j�x�({7�\鑲�������6�Sd���qy���O�t���C�_�!sDx�kyeԋ"�;���QX��N�ѯm�}!d<��&n����iR��d�0V>+�q-��4��1ȼ%�{� J-�o"���\���aH�g�Cz�5s6%�m��]V8��ܶ�-�����`h|A(����4n�`t�V�ǁr��� '�������� l̏�H�閾�o�6^G޿�W�vو�8f�R�W]�e��R]��Kۯ'bR���* qp"`%�S����P7"�J�_�+v�������P����Ϲ� ��/6���l���CT�k��~A���ϖf��+��d�M���0�"��
VB��]c�9�%8��;�Y2t嘭����b�ʍ�>��9��H���~�5��,����ѽ�l^��k=\��8�d�+&c��	HZ�Z7�g/�<'	����9~��獢�y�$#x�/X�.��9�z�5�̖6u��!���t�ө�E[��WYm׎Kvdf�q_0�wB��1o��b�Gy�%]w:��f#�2�<췖L�� =���m�{��1v؍ڳ�o�+���@���|U��#j�4�e:�J팕.�bA��n+(�g�s)�3᎗-��R^r01�\�����Q��f;_�iQ��Ϭ��$�M���"��ֵ�ݣ^���6��u���
��[���XD��}VU��%;�m Q5c���_�q�,�]1�B�" �Gi�C�Sw����S�4򢚍�.�n�S�З��?c	�'�s5��6ߌQ�O�V�d��^;�*}z:�m�T�s�G�*�d8�c�TIlZ�Z�Dz=�3���"JX�IⰅ�^�U�)�.�M� �i����ٵ����l@�	�8�naULmR����TB�����:{�=�b�O�P���h��Ȑ9x�(x+����}]	g-а�������W�.�U��3���9�2˱���~+�&4G��(�T!B� @l��/����)3�_w�������Ec�n�\"�1���U��w|��0o�浈��(o���3^B	�Иb`�>��$2�sk�ꗔ���nٲ'�� �5ʉZ�*���K��v۲��*��~gwf����q$�61P&;���	�VQ�����$m���n&�(�0�y�3<�ɨ-m{5�$Շ����
��,�O���� �w��Xg;VW�%���\����4��ԃ�N��;f�1�q����;��k�伝YD�L�ft,�4�6|�@�z�_��'H�mJs��0R	�'��.(ǽ�A:���1B�W>��*�T��-FR��BG�t����Ú݊�_a$~J�J
xF�B65G���� +9���ڃt/����5^���d����N3�q6̹y8�)� �7`g�b������:�~���n�����(
D����NCd�+�'Pɹf ��T�x��[لQ*�c��mZ�\�_5½��c&�z�)�A�)*1 '�)��U)������f�C�4�D�Z��k����y#��t�N�}��Ϡ�����b�\:]
�)���Hy���5��9uLj.M���0����%ٽ;�o��7�,�xj	|�*��ke�2����w��ʊ�� H�O��5p��N}��b�F=2o�M����jT?*l�H�H��T76�~�� �aۤZ3�I8B��|��P�CM��:n
j�OT�M�2�2����D�\-�8���R��V��6�2�Zg�loL%1~z!v�����6S�)�r���uKw<r�R��y��w�d<��L�.����������ƕ�M6q�=dhM��i�'�NL��:�c�1���F���A/��D����%�/&j�Ĕ���B?�~�M���@e2�ߩzEV�G��V,�hV�S����S���Ү����PX��' A8������ߌP��#��4����W8�wϏ��4��У8I�Ֆ=���5�%wp�~���dS����cG�l�Iz�5�-�A�] ��t_A��$�U�@����	�
�����e"�!4�:��+z�s,�=�eVZ���  ���M���~=)�*!GBxqm�W���,1���E��H�7ˤ�cǧih�2�'#���P �~����2�Z�#n]X��Z	C����ӆ��	��4-�c�R���濛��L�T�@ +�7xs����o{Qى�c���%��ʸ��"�����4���3;��5�/�nU�oV���(���|ۯ��O�;��<͢�������5�z��o���M����Tt��*�,b��啺�5{L7�P-�O�^�&2�G�vG��g�hG���K��~��sO������&�ԡ��3�'p
>���FQ/�7|����h�$
�c��ݫ�e
��Rq.oE�%�I��z7�t=e�����5�>=�ً7��f�=T��"�Ú� =���w��G^S;��A<�QN����P������+�]�啫�J(b�<B��O�fd���
S��M,����o��9�8�����Q�%#0������M��M�ox���a��g=j
�q�����G��8�d�x�F�HPB��W�zWL!���2��=��y:og۩4s�^���zB"���[��k��� 7}�@Sn��P�7�o��iA_���<�v��wmI�����sԛ���ԝ,jUK}��0�ѣ�^�چ�����m��[��}j���Z=<�	�W���+���ɡCב,��5�@���Ɨ���Vf,j�+w�CX�/�n�rV5�b�h$�S1Ņ7A���h�0�)ٿQ��iL&/��&"J�Ǫ9��P/�F��'����0ƌf-�n3�C��Nx�]y�paٲp��mǳ�X.^���2CУ�esK�� ȵ�e�����$S4�IͲ�B�;��;�ю������U2Zz�fa:��fL��:N݋�I�H�����ً��Oh��i�$���cX$�N���0�O-4e��WL��;��"�����;��s}�+�bm؞PC��C�,�a	*���}M0��vw�/�����6�����?�����d�j�l\32�-xQ2���{�CD��o]|gq{���2���@�Q����I�1$y@�n�ь԰���|�llg�?DiZ�-F8�oe�����Uܜî��՝�n.��{yD�9�?����ӏ�]�b<�lU�u��ڕs���/�$U;�Dt�����X�=�/���q��J�ò��Q21Ɨ�ni\,��W��Z1jYTgzzk���P�i]��u���:R�뱸�X�����j�h�+��䋎�2KUp4�s��;�Ǹ�|G����WMk�/�{���F%U;��G�X�u�!�ü��:ÿQ��$4�$� ����0���r����6��45'H�6&S�����f`��헌��ٲ�?�y��`'��4�Ě�M��Ҙ���uN�|��vo_�����d�=�uM�L%��$�a| u�R���
+��<�-�CC�;�N�*�m�Eʙ;�Fy>�FE>y���1]a���
EY����z�0����=�M �ԯ@��,��C���J�L���x�0&kQ��@ן�F� �A$���ҿ>��/-��kcEw<�	�Ds4hq�5Z�PFL���9&<~ n:�p\KS>l�Ĝ葮=ed
<��~9����v��S�_���cڨ�è������k�c:{�*���[�(�"����>�q�����ś����/x͵�,�g�AG4��6S����ˈF�aN�Q}���}Q����@��֎�8b̑v��r���S,���:����������0��pb.�� �pfNuv�n7��y�����ˤtԑ>��lm.�1�칈$y]:2|&b
���rj��Ɉ`��ss�OW}�����:�>A���08�Q�RzCʰ��C�55Y���1��3�?�\�7'X6lqjWzI?�sU��xl�����~Z�����*r���0J��'����rR�V��H��70b6T���6����d����kh{���[���$�BK�F`[;Yt�^�v���5,��]�(��ҁ�2����K9�Mj*.��4��fF��i��"��c,%�[���kşI�����l�9��oΐaM}�l����n�� �Q�1���Z	���j�{�6�f ��bG3r;�p�x��� ����0Tr�|Z3�[��m��qQo`%��mW(�;%-��Y<��"(���s��Q=ȷ�:�$Ǚ�2�%@�����?]�eLl�ʻ�F`%]�j�zI8��J���AlKU۩��~�Jv<��e�\>��y�T���5��G�he��5Om���d/IE�D��c �r�qtO�K�-��Ev�`���2��M��v���)`]��V^`�hy�U���5?ڃ�৒���(��b3�D�ݍ������̳�GXʞ�h���������q�dD�{Vh��q\)#�$��45J�Z��	��L��
�����>2�G�	1x�r�ǣ�KjxP���q�[�n6/����>����c���E7���Rg)�G2�.Kt���1�����+P����b��M��U
b�:1N.����eL8ݛCZ�Lʇ���ɏhǵ� CJ:.v0��{l�D��]o]�y^������K�Aq*˄������ȑ�a�qwi�������
��9@��A�|  �-I^-;�pMxN�ڐ����Ӗ����i���ޕ��-6]/���v���@������1�ǠN�͸A�	�7˛���@����7��V�6Ƴ��C	VM0�6���x�g��/6��G]�-�́,pV���&�a��s�!��&�T���Y(J�H`T����C�Ic]m�t�'*m���_>5��*�Kh����&�L�@hƱ��3n��uXwHH�¤�v�yV��Z�@���M�
���mǳ]�%BE���f9�֢��:��̂il���C����G��t��>�n�'O�_�MƏ~��݃g�:,U,�>�kS?�ʗ���k����NC<d��g~��a4�!����R������;)m�(PQ2)��tT#w�?:���&��w��$�]���q�Ck~	Nz��ct,]l&�ڛ[�%J��g���^��s�Cf4���#�;^��"��u.?L�e��
T�Ms5���Q
��Y�ѓ �P��o��Y�
�j!�j�z3	p=�M;\�C21��ur<#\T�0��#d$h�f���z�^���ۂp��vz�鑼�3�9jn���x�%Mm�s	Pi��j�K0���вk��j�"��A:����g�ߧ��2��Bv��|~���[Ai¶7��4�Tߩ��AY3s���x�>n���;��S�W��l��? ���$��j+VM['q3z6mh���ƚS�d����Q
^,y��A
U��M��hh�x�3���r����	��o���I|�`�ӓ�xW�f��:L�V�3DK1���gӋo�f�ͷ#p�3�8�[�� �����@�*�����f��{�NOc�����Xl)�܅�9Y�P�=#�''i�����f��&�a�^�8D�2v!��?�`{���,$�v��Щ�Ζޖ����(v��U�o�o�(��3���5��>�
� `�X}��O�4RB맲��?�D�(0�)�ft@>`ȫk�zG��d���X��W͵��o`>������J���ae.S��3f��iڴ�a�2��q(��vW�� aES����f�udb!|�Lt��s,�����g ���G`L�ӟ��|�q�,�����Z
�K�_��X?��Y��%30xJi���n���/�����¡0+nf������Iݳ|%����8f��#�C7��f]�q��:bnݽ�£��w���*o"��5 L��\<B9=�؊�����G�;��-O���Y�wJ�%��R�uk���7s���Ĩ&ͽԠ_Im���a��(#JE��]�f�1�r"]��d*���L� H+�SD��Y�m d���R牏	)[��L��6Ŗ}v�ɑStTF����oq`,������As::�oxDk�Ctoƒ�@t�t� �/n�$�����\>�q�Ⱦ�T�
Ȫ��9R`S4 ���Q��^�]�C�邊
0	�?����}�
�>�R��Ư4.�w��~��e�a�X	�'�)ޜ\�*���l�L��|�K�a����h".C��gEs	�QQU�[�]U똴��X7>�X5�.��P�
�`�F���,9?�{P���=�g�p���glM��N���/��r��������HPe&8�醆-m�#I\I0O ת��!Z��+d�d	�kz�g�w���@��=����X��͔�.��ޚ�aV{Cg-���~�a'<�_�!��
�ڐًS���j��a3��"����_���|.w�&�p�[��x�2� �8/$j����4��Oٯ#U8]C2�Ϭ�X�ks~�]�{�g+>&yd��F� ��FD}du�Ms���ő�4��rSI���M���H�rhg<�������qt�dR�zGI1v�!���l}��	���)���ԱfB�'�`@TPRI�|�8�+ GE����W�T��2������f�}e�[�Oߐr��]�oz.1M��s�qM�9V:�Ϳd<���q�)6�M.L�7�\�`�t���N�'�?5�wһ�ij���Z���@={L�y)��ɜ���D���c8���݊ݯ��@��$
R�e��D�F�و�0��ԈƱ�Pʝ� ��`��_�M)GoF%�F�mā���B�^�d���?y-hՕ���8��O�l1�S�|�:%+Ô�^�tZ����*�����5��Y~6�r� q�=�8-�g��Xh�ؽ���uw���=����w�&Ϥj0u�/]m�Z$s���B���zv�I�	\�z�3��>xG��o�IkY
�j)�a�٪a��N��}�����4&M�	hex[��_�tMxJ��Ʉ4U�9���t�p�#��@q�$�$Ó�\�ɤU����#Q��5T�^U5�qnT���;�!g��N�L=��~�ߪɖ���ڛ��ls�����zU�� p��0f�+�|Z:��-���E�b�qD��;���)����0Ƶ�!��@�y����Te�k6H7�cܗxwT�_�x8�5B�G��wd
3�+3�:� �Q!�/ �8����>��N�u��3`��	=��&���@���z#�33y��B�]�:- 3/#�Ro��>x�xC]��i�"#}�I�c��o3~��Ž�$6��J���e�Қ,��͌X�-��V缼j�,=~9�4)O>i����+��f�1�����>K���!S�i���/t�~��?B�䗰���Y�L�� ��hg#m��Z=iq[w��~͋�� ���ϟIV���kvz����n
n&��s��[��6 ��9�H��S�bQb�.WA�D1Վ9���&s�o-	?ws�X��M���m��."U�%W![���a7|���*�Z���� �����&��Q�4�<,o��n�Y(�&�֫V&��A�����tɅy�8bt��NmDz�G�w�.$������/2�Gca�C���i ��%��t�"�������)���]z+�C�I?;"̣Ӆ�� ��)/}�8C�Ba���)*��c��u:7���Rp�g���X��|]{KX}oLG o-wj2v�ƚ��&ʴ��-@iFt�s�k'�{cFmUh�1��m�%�O=�E�tZv�r~a�+����Ac1z���mr�6	̒$d�[�� 滉d�b�H���\��A�䫹�HW�(���'x/���HV�m|�O^{%/:7��V����
D*���>\Q�F�-�sI�Q8�)4$�隍�l�`��Ox��q��@W�����;7x��"��6��F�]v�`�sM����|W�DM��"��ILB�2��.FUY\ׄ��͛�4&w$Ք!�}�L�$��?��$�4�� ��I`��4�K��@İ`8�ۛ�U���=��N�IC����B�7HiY)DoP/k�����o��8of]���C�p2)ofĆ �FLJ֘��ANНy"�+�����ܸ��L�K��&�i	��&�L�B�/�⿨:�!y��b��Y�I���,mZ���u�	 S��3�:\ǷT���8�Z��sZ&ԯ>�̰��N���/-5o�s����c��7�.P+*�^+ʳX�wč�̿X� _�
���a��.�葀���y����bc�R��U����{R�^���{@��V�G��X�@�GB�FS����4=	#3ҶE��
i���SY��= �� ����-���B��`�o����P�T��v�Ѵ�t؀�e���<�t���FҒHV�xN׹��L�&�����e1��돹�΀�,��%W�c-�H]��4��N^�wQd�9�e�8�A��`�g�)��[���t ��7�[E��B�j���pQ\�H���/�ZH^�@8�@t:"�#�w��])A�oږ���*�.ԋq�
�����hZG{�|,�`�kL#Ȏ��6���RpCy��c�yz�������a��Q��S�r��1u���̃D�B���ڟ�oJtFe*�
��/s��>���`��U���AYG�a|�]���Lq�����͕�Zl�'�����n�DP/X��.+�z��*?	�Р�P�wvB�k��u�	�1C8�|/�U�g�;��*Vz1�;���~�I�;
ɹ�Bϴl�C���&�gc;�����rm>J�A��N8�:�x�;���+{�
}6)�
oH�U��-<-�3�|h�';t(B��_X<���Fc��l�]�L脧Y6E��H%ggS�s{pMΉ����2
h̴�m�*i�!I6]]�d��N�@���2E����`��s-�XE�<�^Q����G
���]�3�̐�h��m|W	!=H�j/.-�A�ok�sKq��Ͻ��~�[�����A� ���vxe7�5� ��M-�a��8�)��W:�f����l��}��ߑ��5G-�<Sy�'��%��v�������o�CY4�]��+3�aϬˏ���A�I��6GYLF���1�����rL�p����z���#@#3i��0����i�4�}ZqU@5Q�^��iy0�jd�m��k��-�2��A���4�oQTMUG�)�Ɯ��9C��u�j*N~��/ ݿ#���\'�\s�%;u/��Dp�_=��I��R��;��<l�~�쌎��^�i׬�,�ck� t�kxG����p��g�}t��1��UEPY:�B;x�W7N}���L{��R<�{�����~�);d�·W�	�]��R���
Tۍ,�������nŰ�Uj&����󼃼���^���������B%	��O�IGoD#y���j�3��*�A9�`�BjLY��zӏ�`x4M���aK��Lª�1�vm�S�����S^�����ъ4췈�d�:�?�@�ΟG����>E�50�q�]d�e�?���oV���2.��L��bk���w7��w��eCB49P"댞O��B�2��HcFm�f}Ő�y��X��Q�{���=�������L4(��T�hQ6{�ʨ�j�(R(����ex_<"��>���	6Y�!`h��؄����SSٕ)�U8y�6g�5Q	J��34�q,�7߇#�?5��-A�t�x�B�_��k�;b��b�K�N�8y�I���^{Y�-!�P��`�co�l���e�R�%�*��ny�p���J�	T������"Ͻ�ŷ�O���y��L� �L���tɂ����������zQG�L�h�_��|��W A�=���(�l]�{���~��\�[q�+)y��t,Z9���ڷ�:���������6-��ve0����0<�'�*�o@��+�l�t7�d������yo�cOܐ� KqiL�NF��P��_r�z���pMp�5��3��sۧ�\��*..扆#P���J�~�O�\}1H�ձ���"0��J�'�.�[)����� �+l���X��Ľ0	�,S�mi�b_/�5	��?��7��e�Aq܈��pv�S�F����Z�t�(D�	 y}�&�mx�=j����F3�O@�$o�f��;�<��Ӎ���~f}�p���iȈ�@VP����l:�B�p��99[�,I0��6~tx�������tJ-��:�r��`S�h y�!u�Up�J���1���H�i���?T�x
�a?�n*�`��uie����$,�<,q)P�+�B��~ٺ
���j�x�5JU( ��g!��ଏ�3�J�U7�E?5Z��X�z��fL�XӾ�@]�yX-(T۳o���3A;�%D�tj�/����<n����}5��Cj��eӬ�ڧ���y^�%c�;Y 5�n�����ш���$�>]�`f�:D�c������d�7�9
W�>�G����������ڲ��̮��8��rfը�[�g�<��IufK�&0��G�m��=��Ǔ/�Xc��ӾkIB�]y�0�3��S���&1Z��>܄���B�u靿'�V����C���B���q�;VSF�-���B���KᤘU?�v��{;��s��C4 �U�:�)5#��<��_T(vۢvQT&3אY����h�_��1Ͻ")�7Q��)����m�2�6wQ�햛��Ka��w���Eɇ��x�X�JIe�!v+�M�'�ĉ�23��<�E�[��fѐ􀻾3�`o�e�cԆ��8��s�*Bi�B=C��#�u�j�*H������(v_�FV�U�s����L�O�CM��0O�zt�-��V�k&��"���9�� A�߷��W�޾69\fB�ٰod�r_��f}�=q"Sŉ�i�+����W[Yu8z��j]�{�V�C:U���Q@<*�3s�1��p �D��UM����B�QĆ�ϻ��l�؎i�YUh2��x@�� ��27ee)Z��ƺ0x����q��w�w��֡�P~%M����6N�Ț:^Ĭ�)��;������d�^`��aĭ��qk߱Nn����c��?1u}���:�@1���>�h�;�DY��� -7�)!��`d��GT�$l���P:�p�_S�p�̋�1���j�)`s����gn����h�vNI�X����:��*{x��F����Ǡ�U��27Msa\�WK�(Ѳ�����1ّ9�#�h%�� �D��K�uBE�$����䂜��u넜���������:��V�
�a��'t8/�_�����;5�ud��E�y��bht����!�w��{n]q_Ց�:h��nYΕ�[ۭ@�:no��L��<�������YՆ	�o�x ù�}|A,8���lg�]�(,E14-�K�5��j���{������u&/�h�^�e^�1�X��s�6,x	d.J�Y�rN2}ք��4���ԇ���	�����|(%� J茰֕����>/	G8Fh��I7d�$&f�,B�Ax#m"�`�"�aK.��L��j���	�,*A�hZ���$L�5����	�"P�43/�0 F5��x1"u?�Z������]�ڱSp��|ѓM"�X�Hc�[��5�6O7�:��t��B1�tm�����{I�N���p�
.-g6�c��R��[6w눳k����rS<�ŏ��
X�OQɃ�)�o[Y#��_ �����P�˦�\��,$���7d澨ո͈,:��x;��0�ʧ���|�Ď��쎢�kr���G�p�;hO��	؜���`n䕿DA�L�*���&�rj��Q�b�R��:Q�3�rΘ~�s��iJ���V�����[\klmSݿ<|���j�M�eQN0/B��Kd���3g�;�"����E<{Mw�<=l�_�#�U<����GX+X��DJ�|���I��ܽ$��E�{I���<ܳƙ%��%�LѪ�_����ޣ8�r�����)9�X$�0S��KjI�X�^ڍ��a?H]QD�%M����YEu.��krM�6��g���u�F����pܸ�8/�F��f2w������n5��r�|0dW}>Úb�fV�����Fpw'Z�;2�e��-���G��_��bd�io50oN�u������������~-�����^����{+@�v�������:B̈́B-|na��':" ���ߕ��^b�{������Q2!��Ͽ��X��1Cm�nN'�؁$�_��˸?����I����%Ԑc��$@iN�H`�)j��@_���%�Oq�r�/fraO�~e�jhm)T�$���.��s���c&Jq[c�a�uY���s~V��+�B�}Z7��z��?t��',yV�����՚®j;��Ξr��=�[����\L�y��:�$���@�1�߼��:���#cN��X4x�->SKzY��-&7C��Z�g% �km�TGTށ�PBPw#Z����LO��D��^ x,��-+�W�ēW�8��'+Cb�SMU��v�ȫQԈ�Hi!��z���p#oa$�,�3e�~�v�睯��8��_�㐾���e�J���'Q�巜�8i�.�JʱHJ��l��,p间T׃$4=�k��@V\6n����U�?ƔĂC3�xJo��q�}+���U/@�D��y��E/-��9�d��E���M]����ܠI�Wg���.p˩aM��k��'�t,���"U�ȊR޶�Cnh���_�w�=l\���Þ���=��g���m�t<��@�3��+�m�y�H5�l�{��ud�Ӽ��>��/�g��WHQE�����3�/�����pc�$%)
�[R��N{Hgb�h����(�����Aj��1�7���J/� %��l��,,Fb��,vi}�R�?Hf�>)X���}�(G��ۇy�ÕJ�i=�K{�5�dl�4��y�dK3ë�g_�#�4���t�������־0�+�_n!�e�MED�
��,�5M�l.��7*DX��P��n�'T�-��?y<��k��Ij�<��Y�x�6�CJ{9��!���u����g�I�f^���y����u��o�&�)��wb�P�W���`�x�2a�*� Aq��C6�X����A� �+�	��ς�
�o�k�.�7��j�:��d�:���z��^��	4�+����!=�Vq~��t�x�T%3
� ��w�?�G���@J���<CZ?#�e��]o�[9|���֠�&V<���V+��f2%FG�0����o F�r/Ű��e���di��8&��_~�ms�}�n�M�����'jVݟ�h�W�_���H���џ<N�^��&%L���e=���ŗ�k��d�C;��h�+�%���E&��6.��vy{�oف����#��[��T�n��f��E˸&+ڀ��Рg�M+C����z/�бV�����fD⋿7À�	����ֶ����Lm��Z��^��2�Q۩x_��ySg��S�T�������5Ҝ���8���ozƣ;lC�j�z3 :f^��L�9�B�fؒ���2K��Ƹ��n�g`g����+�:�v������/�H���^����G�xnU�H���<:[pO�*�9sE�@�aOh�u�}V�	�ijSL������.�K�~��	�P����4;T�|kz*����Z��*W�i���H�o["��F�2�y�b�����48�<ɪ��8i�۹Sc�%�E:����#^�ޱ�������s��"��+wס�xSrܣ�޺,0-"pUV����y��'�<�o�I�P�?�g����[�g*�I\r��ˠlQ��"L2����9f��®I�c|.�ǎ�*�j^�P�Z�ݕJ��9>�i����>�o�n����[�t�I�9��Fer�߳"�LH�k�y�a)F	9��k�
��V$R��w�n�9q�����ְ��e=8X�׊˄;��TLJ�Y9k�0��h�����	D���y9���6q|7AZ�b0(P�\>,LMS�QZ	�ol5g�1��[��k�S��
EK��H�+�3�����q!8�7�;�ᲊLO�05B�k�[�'�/]��6����O���0X��!��A�����kayK_�OK��z�� E:�w^�5�SCU�,EŲ1���,��ݹ�<]A�o�T�N�n��.�ف������������
Cy�Ԯk����"xrg�o���GI?+0M����QJ�?PEU��4ᣥ��zJ,��If�ۑ:�7,��ي�ɩv�[-q��V���v0`^K@�w�<;g�%��
��G���پ۱B<Rs"�^,���[��Ѧ�d��U�����ڭ��75�-;� ����X٬&i�Y���Qh#\98�l ܚ�8'u����V�n\vRϓS�n� ���7�HE��3E�.H�-g���CO����k�Bb`J�g8�-���0�(��]n|3�|��my��u	y\����E�b���7�h�����
"qF&FP<uBW���$����ԛX�x���7�2�W��5D��ޚ��Pf.��A��'1�{-mŎ�+�Jȡ[��mˇ�~��㟸�V23}��D��O�-�C���-Ցt�չ��v|��GP&��WM�S8&�6��!�E9�#�P޿q�*��.�����S�����5 iz��w�kC����H.jN6,�N
m����o6@�np>�
%ۑ�r����=	����х<#w54ڋ"y����Z��7=I���*�m+���s�Y�n��o�ƃkL>�ּ�]z$.�e̟�A� ��Z�J�2�\�B�Z4�o�qc0?Z�7�zэp����DW<՝aV���-��4�ㅶI �G5�%�U�ϓ���29�?�j���y�%��t��,{Ar�	�`�~ЊX��K���:�*�K�a���%M��C�ֵ�o˼G>U��t Uɾ�	�(�9���r�r���P֞�H}��oS�޸��ki�ք,)II5e.v�
1v	t���B�R m
GA���E�%c(c~A�G�;��XB�A�>�gL��x���C�t>���wO{��5U].�Q�!��:7Ǒ�M�Z��U6�VOj��.X�2˔�*mI�ρ��É�p^2����W����q#�d �Dw��сT�ͻ�7�(]v��� �#{o��;���^%�JmtQ��AJ� �eI���p�:��$�)�u(ՌM�w����b�l��f]�̑Y� ���W���q��I�k[_L�OC*p�D2o�	�b�����Hн�:cΟ��hz��,:,�X-k|Dn�CCKYL�<�7��F��H�c �bk�q#
�-¹9c?m�Ay�
��=L�Z����Z���
oڑ�C �m5���8����=7"	o�
�����qK�1��ۿ"�V-i�P�Lm�	���w�͞Ww(�,2[%�xuJ,�C��~N��Nt!F;���i��U
��qp��r�<� �1�<�w}�X�ZԤHoJ�1���!5S����f_$����c��p��6�v ��ZcV�"�L�7�Jk�b���;��Ŷ
�yQYL(.<���޻C��z��Xp���j�P��� x!;�˭n%����;�q�>�*T�)��T���g���͵ʞ^f�� ����L�m3>�����^R��[&���:��|�gw�����|�����tt��<��F��P1��]�G|ƅ��՜*�l�p�2�=�d�(^nA�'d���(o�M�9�ERB<!� )��������++�� %�~V&a�����Q����Oa�]�� "p\�������+ �����s�i�����U��̜�'�o՟8���9s���r�D�OÜ�0s�8�����?=����7�/�|��cu��/	A�[5��8�A�w�9��Q)��8C����u#�һ�����b������hdJG��9�3n���l$����ګ��'P��Jִ�������"��2ϩ�(M��H7��ZVn����~e[�2�v1U��͎��`a2�bk7�
����R�o���c!�^�C!�9yw��QC܀#���9iTXX�?��o%�LMF�Ow÷w�I-w��'�����B[l�����x�?�nv=xVux�u~NOl}�|��I���X�4�8����#��?����e��QpP(:,v5 �Ft��OW����7��|r�=C[2��J
f�>%���c~��niۤ�}�m\��KD׾��C)�JqK��ѹ9���ձ~���fk�gþO�J��,xh�u���� ���=#rV>rG
z|1����KG��E�I��B(�ge�}°���1��;����K�� `&�)���k B�m{����6��������n[PbW�y�|�P��:A��Z?� Oe����.��n\>%��d�������4����̆��cAqX�ʅ뼾��T�o7=�j9� ��2O��X��A���Ә�M><b}�<]�+���:�
r�ܴx3e�����ѝ�����=q��Z�����U�p����p��~6��UWY��v��kt>�R��A�]��[�g�񵵗\�M������Sy�Mץ�{��#�����*�����ePN
���<��=)-��Y���Ȼ���%Q��=Y��!/�c�k��HJz6���.�b�|(�B#Dœ����m�����WC�%��e�7�Y���$�}�y��+Ȁ����v���H���}1�wm�g�ѩQ�[>FNq��s�������%]jn�q�W:�$�g]����]b�WG�="�C�d��)�&b�/H�5n�H�LO�U#2�����xL�������D�%��f*���������ی���p���]×�V���9Ѝ��֖���!M����^�`Xƭ@.q�����dn�>��7���G��'���Fon~�>V�x�^��F�d!fd/6�~d�+�J��*���ϟ�2�Og�������� a�:���UN�sX��H=�cc'O7��cCg+���� m����j[#T���;eZ6���@�U�Ŝ����!~�����A
�Y�y���Uu8�s��L?h�E��hw�>��Z�e㇦��~�,pS������Qt�F�l��T<f���TKr
� �M�\��Q:�e��!4v�^�l����I"�6��2�lz�w��u�"5�|����q�eh���Ѣ4^P��߮i�~�f����eCz�!��Y[O�����Gƙn<};2v^��Zl��,-6:�4���HF*5wrN�+��et~�a:��xԒB|���P�FN��IKhG?m�f��f)K���{1�[GI�v	@�rRT@�eqx%�Ä&=7G1��m�H2$����ٍ�:T�?���=��Hg6.z�<���C���K<H��������9��"��+gc����"���YC��]֭,���a71�.�����<[���/C�&���X]W'�D�[���J�T�\T�3�U�~�T��2c~qӊ"����NvD�a�7��\AZ�L������x�?�Gi\����g���'��Kۓ�e�z
z�-��ɐcR٪;��m
+�����|~�\jlh��ԝd���a8�`�����atז�a�fʛq�t���]xM��v %'7���?y�=��c\���u��[Rf�{�3/tT�x~�	������[&�{���lր�\�3}0�)MJ�w����k�%�e��~��1?�
�$����"�����y�I��8b��]�uQX|� ���43*n�ĵ�r��y�0_��t-�?+$�l������I1�X���L'S`*��4�9X�',��\����"Fu��7_<�������H�O��`ܼ�	�2�Y�M�2����oY�z+�Ƶd�"�E��\�	�Q��ƹ_2��������/���`꼀r�@��������m{�s�s��0*��L}8lb㒙[Rn��B�[i
���m���e^���˭R�3[ *��Wj��/��B��I���?�ho�=��'	�r�;׍M�xh����~?�Q�8 n9EE��o��gݘ!�_��� C�(����������{!	ͪ|H(����0����.�ؾ�̭�}4�� ��W��؂��2a�]xӝ������fC��c}OX a+��b�U��9���Y�w)B�B����Tn�rwT<�I[̘�m �b{tvҮ���>�1����K_ߐ#��q�yXsA��Y���k���_�5�|ѺH�s&l+�S�rÑ���Xx�շ�|���r�B ��Jvsr,����c�"��H�A����C�X�C���k���ʔY$A��V�$����`�&]�}��(�F��E�^�d�GJ�V���%�~��Or*����쯾�㵈U��f��L�z�5r+38\��	�BѨ �2�
����	tG����&<��#�Q�q�ߕ&Қ�L.���Q���zdQ8*�C�D�E?��M��v�ɑ&6Y��cyW�]7�/?�V��|6׆�?�*	��d������r�}���{f��7o������gY��crvs��|0�o���ѿeRZ*�#�kb2���G��W����6��ל����G��G�!�Ͳ�[\�h��0�g��1M��~5tR��V���z� �8��J�Z��U.8����>7P�� �.<,a0���p����
�S��XKR���1&��k0P7:6���Ǝ��.�f��g�/n���A�����������SRj�ף��Ls��d�m�0F4i��N�s)T��,Ӯ�������V)x�)i�V�)����1����-��_ŏ�����"��ī�Ǣ;p��-W[O�O(4�k
�RԇWb���ӣA0w<XډeQ��	g��L��FM����ⵢ���K�ca�p�]��iO9�~��̱`esH	I@�-v�vG�������������2�'��i�!	�bdNkz�k�rz��R�=��yB>�3��`:#�zDh]�892��qRF'��Yʇ��:}%֘���T���������Ѻ.�(8}��/�M�����jFgݲ�pB*�q<\�J��LMD��������LO��VЉ�֦�9�q�O:�ȑPJ&�ͥ�+M�qH �kq�s��Z�
 .c��Y��.�U��V�ڊ2��	�3%I��e���g���cH�v��j��r�g�`DAAޠN�b@tRNy��M�� -u1��T^�6�f�9��",F�,��Uց���~K`��	�7���w��?��U����֟�|�To�,_6©�|מ\�����5\*�̚�G�!���p�.&����B9D(��Fזaj����6�7ѕ#�>�Ϙ��[�P%���G�����J��t�&�Wֵ�R?w/��F@�Vv&��� ��~�����l��_��?��� x���M���Y%�!�㳐���u_�łƃI�{1""�>~�[L�00A�&W�T�5`t\���$/5)���+aGs���}��%�oW2��0�=��Z<�ovH����?)4,��]�T��$��\������O�.�^���^x$;��v���9�����M�Z�>jV۔���M��y�����������!S�)��'�:i�(ޮ�^�� ���BU�p
���uf��R�xUH��v��@������؎�cq�2���A!��!A_4�����`*��ua"�d�eR�~��Q��[]��cp�_3�z_r[��o���x�oX�{p�_1b��%S��yˬ�$`�5MV8$�Vi�EI�4�O/�9��!��|�8 ]�.�W�h�o���A�L��u�@+����H#v:;0ܭ�&�~�@+@s�Gn��%M7J��J��8�h�V%$��B#jP-)Gg�P���(Q����`��q1�Ii���qNmuC��N�
}��l?�@J���.��Œ�iO��V���ym��sCƛ����Ca���yCCn��E[=��x�9'l��C%���O=���<iS}������f�gHlr��2{Nخ?�-��o}ER5���߈�#$ۇ�֩c�l�$?0\ak��.��ն���n��6Ѳ�pF�?��|	I�)���*�m��
�-�%,���.��u/��ej�J��ʭ���������H���}��nO��z�1'"b����*�E5g�IoS�Q,$�����=���bAD�� >U�^��Lu�]#��By��	�:�3�qd���u�T��\��dE��*��%����sb-Ј�=C�LU2QQ��3"�K2��8{�[o����)�G�m�8�z�(Wл0n����Ԡ&\�v;Yӝ��_N���f�yM]������a��Y��{--�*���t��X�YS���� +�S��ť���\�Aݫ�AL��zx!Z��ʅ��@;f���E��L6%���SC��Ac�J�]E�)G�A�md��r�2UKAiu��-ڲ��G���t�6�&�о��������C+ �kbn͏� =��u�q��ήy�����Ժ�vP��A�Q�w�+;`��' H��X޾�$ZH��uTT�nǮ��P�r��m=p�b�`T{����k��8;��%����D�*t+�+K����p����z�Ґ=ڢ�h{��X��
p��Ǜ�3�;����J�@���u���F�랄+۸~��%�0�$��,�-�ʚ�b:jZ�E9  Ki���Kb1/�%�T�u��XE'P~��U���+�v���;N{]65#9}� ����f벹�%���u#rB�U�M.���=	��O��j�\��8i��_��q�\�}g�/��4;`~.��.���OU���2���BE�ru��m���Cz%Ŕҿf"(�d���D)P��n���j7��밨g�3,Ϩ�u�����c�g�Jo��2��l*�y1���v&Ð4�bK�
��}+�Gpy���Vj$ʹ��D���e�p?�r��+ߕ���U�,�&v��v ��E�I��CDy�j�ւk`�,��L�Ͳ�/փ�T�q�No~q�s��L�(��ؽ����KKG��hM1\5�*�LP]��I���2r��Xr�
Cb�����B�}��	ϾJo���=�������om0��
'`����oϗw힍��Yf��r<�-R��t��O���6�Y5�b�N����l�Ɠ�����i���i���,���ϊc�H���7����V���D�'��@z�����6A��)nYq�\$���+h��d�`�x��]�00�� `�J��S������S�T��A��&eÚ�e���U�,J�XXDls}{<�y;$�A�;T�������t0���FU��q����AE�K�vLd����.��%ȹ�C�8TR3hͪ9�p���N~�zm)�%"���7��5�2��%�v�^�hHG����	�,�+B����n�f�[ &����}`�(f=��:7�P�8�����X���ӕW�ڛ$��Y������O'SÜ��� ����"2�2_�E��_Y�w���A�TWє���w�D���+�����a�O��R�����Q�)���a=�Htl�;���a���;�HB��ʫ���!�IXyi�W;����G-��!D���"9V5���$�=�p�x;�}��b�I��fX�
>��i|i7�^*Kl�ѣےt@�8F�$CB)����K� ئ[B���f��i=�E1�ky������_������{'�
�Q�np���ꚝ7(��u��v��l����5�}Rl���c�.X0�2l�8��!�Hg�{�`��Y��k�V�J� �F�̬���<r=��9����z���'J�Ma��pm
1϶g��:J�dP�$>\�-Ͳ%�.-k-U��b�rL�ʅ�MKO�IW^SC�z_B�!�ޮ�c��0��)/��;KP`�"+�;!��Ϻ�����5�@IŌJ���CK���[��y��Fy�Y��3���=���$�9������
�� �m��w(C�������W��|��;�w[e	�r~F���Z@�������_>����*ZF����'h ����d4	ݪ���js{:^5��n!�-8��j��`��>H:dݤcW�I���#:�P�
���K����	`��M{��I�N���.�w2P*��\�*E��a�Y�m�R`OX+��>!�͚ꯐ�4!s��qĢ\`<.ma�W]秐VU&�ǵp��N!�O��w�u����0R�8R{�X�����u��(�~���b����SX�J|��=}���<���@;1��Yn�r]S�r��qH�E��9ƳF]�|E��|oW�;l6+Ve�S�f��!�w�k�˪z#
jj/�O���a�#�uU3T=3��da�!���>8�5�uN���i��g��l!}u���'F���7*���,�&}B��`�3$�R�+���I�qʡ�8��L����pI�S�w����|��eh�ǐ�[�6@�t�]�.��a,��؛��eJ�滩��������ax��:�X:F����`=2V34�uH�x��_��j�����=��@QyR!Q2w����.���kNt�$q#]�����W#���\�5���ס��pc�28^˯���r �"����Φ��%2�^9ϑ��l����\��U�WP�̖��̨�(/���R*��o������B��+��[�)㙦��%	�������ֆ�Ҳ?#�-���/!Z'/�0�i�p�I����c�KW��0�E)}s�"�y���� 'l͵�5]�@=�ޣ9pX�>�/M]��YRN�=�����чB*�Z�X`�u�Q�H�P$T|Q�[N��t��dk�S.zַ��������L�*������\��0�\|����|���#���N�K�9�6�b��������0cS��"kG��"7��f&+Y�vX̗`d:�%�ͲJHl� P"�z��暹�M�g@���fjpz0}ָN��Aj=�B�{2��!�N�bmJ�M��}a��L_	�!�oʿ���8��7�BC�Ui�n��0���F���ڷ���\�O�ސЋI�T���l
��`B�����/z�r	W�е;Sa�N�0I,���#ҁ��e�a	wz"�~���w�3����h(*��`�ihS�X}�}��,z�AD 0���Ҏ��� �����y�]`^�� �l�8�8?H�z`V��Q� v�e9��^��b]5�@�e_��*�0�Lt��� "��`�f�q:9ņ6��"�g	tC�ˊ~�<�1�mA},U������������T4��}`}�`u�	+��{|E(9
Y����Ԩ�m�����Z�����Z��ؿ;�.:�Ѥ�0K9ՙ�)��$�h��Б�P����6�a������Mx���|b��.`�Z�ƴ4A�Ew�R�t��j������A�_V�q����b��(��Tg�����we��.�RY��ћg���x�V�4�0��,����K�Oxر��P<��>��v��"�/Vɑ�R*1��;��-0?�lg֠�ǐ(q��q*�&��~+�5B�01*JpN���FS�$�6w�:��`��DMށve��;�,͢��+����o槒'Mt5�'J"-'(UY܏!|�n����>�cA�<%��¹y�3���f*'�d:��jES�B"�NPnUb����Ԩ-8"��|�A��*d:�z$PR߾ָl�)!���N@�W +5�u�d?�w��M���-(�|[���`����H5Wa�C�'6����Pcv�Ő%i!��%�@v�f�gp�T6e�w0�|<]Z���P�UC��[�{��Z]U9B�mh�N|C�\G\�"M�7��R�"S�o/�2�\3����t�i0S$T�Qm4�<?@"c�ҫ�e�ls�Sfb���Ճl�Kij�x�	��%Z�K����.�c���֟K�i�T��e���-���\�T�av���b'Ŀ���4�PJ�)Pţ��a@�y._����)�����a\s�o�����t��{��xT�o-���7�r�Є�0�s���~X�K��s��Txb��O�HB�B��5���G�
#�D춠��A#�Ʉ������@�q�#~��VPS�]n��<#;i�ٌTwv�����>g�{K�of�9�,����/��Tܣ��������L��,�s^]���wN�*Z\���!o��/�:xk�^G�k���Y��Z��� v��ۏ���(�'&B)��w���j�)s��eI���f%}�{*@�o�ǘ�y���j&�3�2<�pt�O�}Q����NQ���(w�oX[�?�����
5L�%��&��������U�/�����L�XU�O���!�S�\;}�$��	�rs8d�!U,.2��i��qk�u�!b�K ���j�����ƶطhB0��d�~#�N��E^P2H�ƛ����2����j�?�BC��c3]sF ���@�ch!���=�W�ӑ�����:$\��U�_fE��?}�S�}˓}���n���� ճ� �!��u����=D��sV?��+H��J�|��xү�����1_���7����$ݭ�PSM��wt*��qM���}s�W��S��!9�C��S�~�D]:[�[_U�>o%,�Ġ��u��Z���<bt�/�Ł�k�)5d]/pV��a�yu�LU+b���4��� ���=6F���=~�����p#iӸ�p*���j\����j�J� �{[(�L hx�Z��\�7�陹�]��[3'�q�*Z�<���\�U�D�a�K��	,%�2Ynq����B[�l��{�z����d�2���kq B�(]�x��)s�7�wn�͉g�팰\�*`#�,���y�8N�{[J�S���P��e��Tk���wI�?؊����*H�{�G��ܚ
&F�!����n�B�$v��Q:��Q
�:@�4<��ۮV,,PrC��H*ov	W
~���|��:dI�k�=�r5���}{��o������L���gW�??�Bn���UH���*|�`O��ww�/����AdyL�X��2� E0�\m�n�ī�+.J��:6�� -=EEE�~����u!�r�a��Z�t�L��}�~���oCm�'��]z�w�X����
y���F�!eqI@H�j��;Ti����,䪪���|�M6�j<T`��m29�.��ZpL)7_ �Q;:���~~7O�^�#�]_����u,V_�=R�*�.Ay��JO�W7��>�=c��4V9^JPDj<,�Z��;Z���	������L9x�͑v�l���sP�"�����	��a"�'���£N�$��H��U�6�Eˈ2oC`�X S.���=�y�w�e���?�FY�����Zq�H��>@R��A����ɚ�����R����%�@�+~.g)&0X����&�J�/:��z�u%1�D���Nm�T~���:R3A�4�/Q+t�
#�]�!U�g�V�lI����������;~ρ�@g��a�Q<����C�C��~y���/�c��2�������o�b��P>�@���2�{�9�/p�!�`�	p��,-�H�}Ւ�8�����1�$ؙ���T%��,:n�ų����G��$���K���\������j�Aȴе]�7��F�{ ݧ����@�c�=�0��	)��X��6�̬�/%�V��e3�Ng\� ���sNto,Cٳ[��5�i����a(�mR^����#2��U�<R*8�	��}}4"Q�R�"��󙒮���o+�vDޠ\�"F�����i��k{og�PZG��&$O[}� �{4�9�2�����qt�o��8�jv��/��o�9>躡�!~@��϶x�)����P�.��D��5�,{2�������S_./w�"���JV�"u�k�A��Rw�`�	���C��I�P�F��[b��w@���H�з�����I��m&�^��`{=��C??Ş���Y���(]-���h�;U�F�v�c�C��X�d�p/�o���
�ƺ�
"��`�Sd��,��
AS�"�Y/�(���U >$�מ�[�j��Y��:I~A������]�%n�G=J�g�+\�W<�X��Yk�K[\���	���u_joH� �����`Mt51��<K���o�8
�O3 �ƙ� �ٞ9�rW��{��{�{?�0��=є���������C�7�ޭ���l�K�V�Z����F��	|*�k7��]�����4\��&�é���+��n�S�D����O�۬��ܙ�������2/��V��d׮HG{�sk�X+��n"|l�!�����l �p�ʘ6��x�'B���Rm��f^<;R�01��z�wEp��t%!�fℒ�|���$��CIC�0k%]�M<�j~���h3^�k(vR�~���Y��	{q~Vɉ́�"� �-����O�{e �A]2�OI���c�u]����~��;��t���_����h��z���N��Ө�?rq����[�8��Kg�i�5�jc|���Js���{��[�����h�� ����T>�Fl��8��Ŏ����'������T�p�O�5ε���%�������`���O�h�k�usrmL]?��W�-"�Y�?�@~UWM��wS�S��W:vFj�a��ҽ��$�)�����F�h�Ш����<d�zl�ef�(DRNw7?��z�`:��7"�Zqg1�|)��ȿ|7�Y��B����*�fiy��hg�`�Y��:_|���ܭ��CR�4�[��f�ߝ��	�+����q�;]M���24mD� l@���e�X����79})S�;�2eHm�����W{1BN�;�����`	�B<��r[P��/K��L����Լ�T]��^L�
���Zo4F�YU�EZ-�$RSj ��K+v����~����S�İ�������W�R���S�:x���r=VS�)�e��~���Ε����?� ꌦ���\�(g��]�Y��Jƚ������a_��!`����[!�z�:VҪ
��y$\�2������wl0�Sa�v��@�g*#;�O���DB���:Wػ�������]�H�?G�^0���0#ʰ9}>�i&PM8�vե�|��B��=�y
+'Q�q�L��@u�]�V%�rQ�90�m�}�-��p��gHҷ�����4e��K�RyT�f����Ĝ �E�T՟9�90�`j���}_�����A�X{���^n��Q oOR,HÕ]0�]�����]t�B��2�G��j-r�������<�pwL�;8t�X�������~F�R���_,�;�ܬ����m��Zh���ݲ5���J��C�0�ld�M�c�<��x��G���hK�͠��Gt��Du�qo�Դ��m�ym�rxi����}�䅕�������W���q/"І�9�?��&��$V�`0S/��4��>f�X� 0��@%��3���Ե���3׋7*���ec>Q�眦D���ռ	�n5:�w�w�ŖK!m� �#�[�/��iᯐ1�1��`���T�u�Zwozˋ���n��m�Ȅ���!U;��b��N(Y�C;�p��mb���.���F W���,�ʬ���A���U�>�?���$A��П-0������K9����/�u��s�3E6'����t�K 
�,Ҥ,N���c�Ĭ�u*�ѓ0�!�gu�1����**��Z2`��8�6-Ln]C���!0� ��[=��E��U��6!ch�w/Ԓ&�Z��%fd�V�ܲ������/BeIM<	^;�)I_قZ E:S~�;�Jm�4/����08@��n��hT�$%)������O�F��Q2b�v4�ढ़�J	HH�Y��M@�}�!�T)c�k�����0�e{�HA*�M`�B��<Þ��X�2{�&!{JX�#��+7�ۊ�U,}���Z��20�u��G�Hy_�[��Sl2�R�*�9������d�q��_<Ό�0>��"�����!���u
]��(xm�e�ӥ�n����p��H�g ������H�w��l��Q���u4�-&څ�v|~��Yj���E�i��7�=��>?������%������+0]f1�*��1w�5g��[�؁&j�[�z������#V� ���;��k�}˭�;�RC�7�-'��*���;�oWݘ���f`0��/�z��go�3|�W/��J*��%B�5���45n���K�MhTo4q$�w2��20qa�ܜ�-$��ldGn5,68�N��	L7qntaiVaR����:�Ht1���.�����0r[���kڶ�@ �C��u���'������������������ؘ�b�����%��a�#��E��qǅu��׵��J�*/NmN�Z���n���	:H9s>-�D��!���6j�iI��wN�m�2ܿ�;����y&�U��{n���
sn�N���	�Ǔ1�������*=d���e������c|����u=�)�è�:��s�?Ӡ�~� V9+�
�uv��q*�.�i�+��ѭ�� N��YK�r�ۖ�V�� �tb+��'�m�2���τ@��cZX�RrHu��N��`S����5Z��;�7��q��MH� t;@<��͚M�=M�z��?����E��<SI1_Q��8HK����S�� �z,y��$���$y
����C��7�h��/� �U<&�$�y�����E)�"��_�o!�5�T�f��������I��'$�W�p�˿��f��/�蝎T�A��T+�>���w�`�4��.�B� U7�ɂ�6ªC+}���J�]�!G��:��'1H¯]�3g8�B�22�fi�"ܳ9�<t���3�`�B�d��2�1�C�X�����I�E:]������p<ӦW�L�a��Q2��b�*��l\�(R�U^�r�Şr
���\8��3�78��ōRP�O��������虝�a�ɷ���6�+P�ySZ�,��$��
p����I�F�N�IK/y��@�
/���.	��%i����4g���Zk���[�t���\����zH��Bs���%�5�8b�`�8X�T<�JͅDZS��H*�ڡ�7��!����C�S�f�U5���(��F�ɼ|��1�k�$���ؾMü`�W`�%�q��-4��o�˔�|�6���ؙ|��<�;*?�S�3K��)#���4c�YR���y�?x^�}�� {��0�_t
��oרJ�(�A�Z�߉a9co�3)T�>4���h~�$�w�5Y�6?5f�������?뎾��	�_��7�����8�j��ݽ��u����a�,Ye�a���G�� %��P��k�D||>.���8F�S3l'lo�fM�9���TZw�AY�X�������w-����@���#�{�R���
�Z�g� ө�Ǚ�t��=��y� �u~��=^|���)]��!���
��Z).�EY:Y\���Ka� "�NE��t�N@ �u��M?��(\�s����� ���[n��G�ף����T�/�ǧ��,�J0/��[���!��/9��+�Mz_oa�:�$���6ʧ|R4��yO�bZ��R��,�/͍4�L��i��uw4}���}3ѠO���̞�b�r����<G����>�3�6�-rB}}d)�����Zt|�������ύXJ�ֻʍW�ڲ��E"��p��5�q?
v��Ia$�a �
T���v�&�P
)X���x���0D��hf���{�a�dpNU��0kM���D�w�
��҇oW^���R9C���@�p�x������1Ժ�Y$(��}�Ν�]��Mc۟aӌ���ҫaۨy\`[[J���<'�P=>sj���X��#�l�F�>��]���ܫw�a��~]s\?��2\q�z�Q��_)?�/�n��"��Ƃ��~nuͪ7�^�]��m��NB��zkPvd��y���誎yz��Mp�Ʌ{���+��/���W _KPr��2 xqdm	��"�-���NI��3�(�`(q�T�\d��8F���Ư����͘E7H�u*�������`ej��t�ڨ4;�Ej�� ou���pƈ�y���A?��1#�����\��[�h��p0���Mx�:K�.`sc(�z,�����S�0uu^Q����[�.�r@-��ܙaV��ݍ'ƽ��=�+Xa%?�V�t⌃ӣ���8����[ �&ꚙ �?4�,�4��H�B4�;Nd)9��ǟ�G�
P�1`����̘>�I�,n~N|?CKn4��ImC�����o���it`*�N_������f��,�@�佞Ѽӛxq��f3����K���$#��K,3	�>�b��K�8�E�Q�\��4�ɾ��˄Xn������_H�*�v���w���5k�f����>A�\�&���ZLA�]ۦ���*n�|�1Q�ﵹe�uwZ���y��B��N�S�`Vo�G	����)52Dz��bd1�7@��m� ����W����؛����2U��8�"������8A ��~��g&�Av���c�M� ޕ�[��q��d<�#��".�д�Ҏ�CѯM���H��oGQ��z�o�{�~�2�L�Q�W+æ]^�h�umX�G�)��p?񛯭���F��ڜڦl��r�tK�Q�q�g��Ko]��r#0��+�Cp��PgV��������͈'h�K:Y�֑�
Ϋ�ƶ/���3>�m�Wp8������۠N"�ȫ�$��xOE�F0Ju��}<&o�l1f+�J�,��H��Ċ��rҊ囕TM��
v��֏��QN �ք��N��.ͪ���L���̝)�ǈ���4\y�>�йx]���QZ�9~�C�;�Ҿ�D�%��w9�@�C�u�M����5l	r~6	2���VH�hu��šp�<�o;���Br�@�D�������;Ha96�X˺�h?��F�4���9x��z�r� ��s�zӄC6)</�����I�؍di��s=Pt�-r0ǂ�0#�sr���/EQ�m�L���n��3.RQa�7�M��O[�/�|2[G͔ky��;�f�u��͆®tz��ņ�?������'�(����uj����y�)�Q��������[]v����P?�a��}/�(��׏!����Kv�j��i���Ʌ�^�bSD��)��|Ƕ�����放ρ��o�6Q�ծ����%H�v�pw�6��Z|�͆q]iz�m�]�~k-����/�;HӢ����
cS�
,�(+\7t)�q�p�̺Hо��w�GF�)�֬����Y��Na��Ľ��$�,�ެ1�/�)o�C��eݱ`e��េV��O�F;C+/^W��R�����w�~�%ǃ����obm���]�4��ۺ�wl���D�s�W<�E��5�^ڬ��֥>R/����}��)wZ���Y"�(��A$��Z�$)|f�sL)ΰ����M���©d�qZ	X8�q�6���mK~S+�ܮ^&�
�q�EA�R�:¥�B䨒�v�FR� D+��m)��g�9U��cM��x��X[@RvD0Y��_rʹ���9��e����>��r���1���m��Gw������e䷺c��MP�Xu�g�?"����Cgl��e��(s�ʫ��c1��g�`{��)���I@M[�-���WG�ڟ`S']N*v;h������2��'������������레�$��+Ex�|Q]���rf&.��+V�͝˶6��'�z�ۖ��xz��_>����ܵ���Ϝ=���?I����O5���T��_;�7l�`�����1��D�t��#<��̤�����_y�ݵ�����`&S���j�3�k�ܱ �k[���4�[�M�|/%_ܛ����n\�`y�xv/�*k��u
��,uя{�/��a��J������I���B �F ��Op]?�&���{&x2��*V\���H��((�������u��P�"��&\��N��v���|H�X��q�S'&��u%S��H�)�5��_}���hP�,�SZ0$�п��ٽЖ�e���2p}�G
�$�(V]&�,�\��^�J��J����@C~Pt�U4i��{�Ň�Y�ƶ�)C�3 ѮYJap��<Ȧ��L�*���s�o�Y��#Ԅ�:�R��)�9�8<����7|�k�F��-e`Yh����i�,�-�{�Vp'�.>�d��������v�(�ߝ`皚!�q)-1�'�e��Z��y�\�1Ϋh:I��c�^~C��<��3���2n��&N� p�"�ˍvg��^~��
Eu��#K���D��Ȭq/o��z�2<ed�'�ZCn3O���i�[*�v+f���"��⎯�W�oԂ\�-�bj�+d�$�WÖ��C9r��:��Ki��S�i��!��e�I2��;Ė�u���@E�.em ��vh��&�/�J���5��N�,H����)kr7�-I@4d�/�1�����Zb��`����1/������M���k�::�"/�*����@�v��{��:�jF6�Y8� �Q��=×p�%Gy�B/�ێ���{��{Z<6��㌨���¯m.��w�Xi�:FK�5�% �Y@��!���64Z�W��5p��3oыnϴ�r��*$'1�UaH�B���^��a(��{y[�@)�Т"~�l#�d]�6���O:��-ϊ�<k��|=d,�=��D}�i޻K� �̣�_!?�k�|pG�~ 5M�vE����#�̅�cnt6��t��s��OG$���[ۄ���|��ƺ�z] � Y�!�ۉ�T�:�i�@F���0�H��񖻭�F�7�'�-��m@�3.��d��8�&�D�r�Z���8k�f0���9�&���(�eǜ�O�嶑��������+X�����&�ph�^+���]���f���m��#JP׵Pc��VWy�<�C��s�5�߃#[$"Apyo����W�������=��0O����fQ.`X&蕨��j�j�m�b�;�4����,<��W�A�r!�G?; w!"� x��޶����@S�O��d�W������j���Uv�T�j��/�B-��ޥ֡{+P<�0��:�Ⱦ ����7' �A&�^*��*D�xo���<�,��w���R$~����4����x�4���2k�0��ϒ(�>�:V�lJqغ�]4b�2�g�h�<I+�W �v
[w��U�HMQb���|6@�4��Z�O��P�����is�[�Z����~����a.t%KP�ocƩ0b���� �90T�:���;�߿g��7��7��Yȟ!/ciSK���4N�ⷲ!q5�y�lp�^x��c�h�ˊ΄L�7yY����XRc�� �j_VC��6��CY�O5"yW�ֳ�?�6�z�4Ɲ�!�Ը�"G&U��_\���L���ى�
4k�$�� վV�#k�Ds��C���uh��Jp�5r�������\C�r[W�W��%ǖk�|L����?uyX����k�x`�����&�U�\�(�! �Y�+5�!�ͩv���<q�@�����q8TO$�Z>�K�������k��-���;��*�`�\��Ms)��ܘ%?G�U�W�����w".��
Ԫ`�V�X�m��lu�YQD�_+�t[�� ٵ� ��Ő��/��v�a\ �V�_]�p�eS7#��웋{�4�7���|2����-oXPՐQ��� �Ҋ{^U��N�$��2�`-:j^���c�JP-	^���~T�<{R������;��i���eg��q_ע	��jI�zYR(��z�A:�
����"u��M.�fY�;�B�K���9t�h�N�%��s����|�=���?7Y�>����?�@�A]%܏3��L
��a1�)��4O��4Y�I"�"�I�GCqV,�}f��b�o;����Շ]�\��u�F0"�	��4�����:/�
����	(k9�X�AS8��|}^M�тpf<O0a<���U���O��=p��g3���k��-�b9w�?|}��&$����rô���΀���U��`E��޼Z��%49&)��π�C��o*	�\���J�� �xfJNA�ͬ�Wt�P��yV/�r����P�]���].�S�XZ�]���vj�ড়�2>�:z.���7��F!�-��X��N�0��k���1���vd���!h�W�nVg�����wի=��8��;[O�,\�ς�A��eG7�l85H�,��g��k��Ȗ8R�+~ۡ��J���Y�Պ��z'JZ�EN�J��zhe�=�X-8E^�k�}GS��2黛)_�����<�O"Hw��~�%8
�R�;!��|�HS#�1=�L�m$
�r)|,�?(���xi�Ս$�<<u���,Uq��S����m��������%��G:�sm'%]y�^'x�v/;��|��&�V�I�=�M�s��\U����;��8ǞA{N���=끎տ��A���/�~�[�p��^�� �:���>�i�'�oY�c.�zɋ�p'՚��3�iUt�i�u?4L;e*Fⴼ����A��n�����<���˶��@zN�@9I��p��Y�T��!u�d)_��!���h��6�=��I�3,e���W�syrU��:��]Gd# ������Y����Hz��`�iOEc������a�dL�f�ؼbg
�W�q����/M��dzu��.pM~��kVW�zz���S&\��@4!]&��(�������7<�F�c������ �`����y+u�.1s��e���v$��;J�|�"B�a6�:�Vz� h��8��d��@�N�#4�5O��H��2�=�N\�dg�ux�?��q%k����B�Jph�Rh�������DK���0�ಝ�kM BnQ� ,��{�}�Z��Um;;>��!ွ������K \�q�����~/K��N��T6�a�KZ!Tw�j�����2�+���ȶ!܄+f�`��a�˂!�U6^J�a�f!��Hȉ�X��eGt��l�VK�!���i�\حM@�N��-��2�Yug��H�����m�&���c�h�"�&Y�yo$�*�ɱC��/��B�\�J�Ә�UeV�o���6��S%�yڗ\mtl��Eg�L�&��J]B��d��Y���kG(�q��!P$@ڠ0���F�ق�
'��C�ĔoF?W~_K$�TY�Y�(x)�`�	�r[
d��Kͨqn�闲8��A��pN�w��~!�e���nVrU{�[/�ɪ�����m���a���p���

N)�>]`u����A��-�A\���xG�(1�I�>��>(c�K��¼ĈW�3�~�®�C�ɺ�~+��Xf^R�����{y�{�,�Y[�@��F�P���\��4��o�ӻQ���,9��z�)vm��;�2�b֦d��P �B��Vc{`kE�/���VxxK}�sj}P��1eN�s�]w�R�yGL��NĊ(D��V���E�P� ��J��v�F�ps�t�����V��*TBE`dxZ(��sh�*3e�#�Ie����{]`h���ڞ1��~NM}�]'�5�0Ҋ�t�Y�<��2A����(Ҧ�<pbLD��Np^�b�[�K��[�`&!�;���I� 㫸�@�8��$�D1�XO��8�I���	�_��A+M����I�.P���VGmk����ja$ &P�]W�1�R��a(��J��
5��Q����e/x��[��c)2՜���:&��gܾ��L���2��f������y���<S6d*�X��]t���X�V��?��=� u�l�,�9�|>�;���}��+W��������fr�L�G4.zDi�FS!�7�&dʕcڨ�ri-q�ӄL�/�M��V���『=��5DSX�wG򞝖ya����P��秹����Q�^<��^�Ŋ��y:�ed�:P�/�l�)��Rp��;����F �m M�9�}�K��H�+�sl�J՝A����Q��h�(#H�1GK����GT��H��k������(����R�����h���4���@�;���1��N������v/�x9�(�]�>E˭����(��a��o7��l���F����j�}�I^�� +7���V�"?��C�W����!t��ΐj~��&��r$h��`K^5��@��b �z��p%�#�t��(��6��\>�������U�q�%6��R�z�ί�X.�5>����>��>��J ԧh�����-HI�C�
��&�?lK@��v��~0�r��7c�̀"v�n��q2M�M ���X"0�q��5��w����-��~�P헭�����U���C��FZ�"����,$�n�/��l�'�a�L�����o�V��2���0�.�����l��-"%�r���R���^=DuǇ�΁�!���֑V��O�Q���y'G��"���o\?�������C�6"X���8�D�I ��~��~އ
���8�L�9�* �.V8|�Q������5ưOxd�1u��\�� ������3���a�IU�+v���QT,3~_��m��1�q{+���2K�e!��f"o�{V6�uۈ��h�u�!��f��`c� !a�4����1Xck��Pę��u����	���ӌ�ކ-rX�Ԫ{ob�� �lzr�~��
5���I�w�ڏ�t���a��No��*+�������u��YV��`@C�9(��',������Q���A�3�0��G�y����p͸6����� D;��fB�
|n���MH������i��?O+H[-�r�;����F7L������{�C��&S��ꍤ-/�L�:��9�+����Ί��N����=�2�T��� u�U�y���S1i�CQ\�|�� @��Zj�@͖�3m��\7G�GZ���C�b,��T����4�3�
O7a�m�!��r�J����+~V��Nmߠ�<�A$��:����O�,�.�boĦO�NQ�v	��:y~8���4�r�q������ƋQH�-0�nhQ�x�1���jŢ�;m�{��1���f�P�"ٔ������o����+:���S�#�g�c�״��x, N!�����"̘3�i�2'�*Q�y�N���"/H�/��1?ct�.���z��Q�_�=�ٞ6�M�w�uØ��wTIڈ�p�PU�b�5[�B��.'��v���ȄN�9�}���m��hQ��W�$���<�P����_��2m��
*�KA��F1z�%ۓ�ڣN�,a~�}Q��MLF?�9v�͜f �+��%	͛�����_�Zm>�<�)�LB��7H����!����C�1j����@A���u��o���wl{���'ӫn� Ԩ=�ȳ���8��FA�_Y�t�5�x���C�7��և�at�/h=�3���w}fv+��i�mSм�V2�-���>x^8kn�ν9����5�I�D����E�ݏ��la�KX ��"7��m�kz ���s��@�X[UT�;G�,��Sh�[� 0 ��0�8n(��*�Rɨw���������~�@Q-�1�Q�]O�$]\e-��]� {8�eT���nt^�G��4��܈�f�B�9��E �#���bWEeJ�5���%���҅����,D�`�w�8�smWGi�Ku���cmf���K�@�ugݭ�Y��-OLO�Q�����B���~�n8#�ŋ[/�n$�=�.��
��FJ\,/��<]#H2�!A7������l?|�\;̗�[��c��d��3)G��$�)$�x�`��iG�K�a��϶��y&����6'�'�HJ���mљ��3��ED�fqsH�gʨ��N��tL�_�ܵ�F�P5���9���fm�b/�?������L9R\��OoG�5W���o�H��.�P�k��|ab.�:�`R��H6�78ц_�?x*�z�/r^[��Ռ��q�ҶL�g3��MiO�;n!��ζ�n��3�Y��ub0D��wY!=u����v��n	T4"��1��$We�{yۏK�ޘ�i����*}�w���}��Շ�M���?��mp����?9'ݪ*"T�����ӱ��z�u-����F��v/�!wG�	�\������~>��k�5��P�$~�$v��>A%1	���J�vpN5��,^E������XEg>�@�T���������b��Ƒ0^yx��o.>'Ndz�*Z��0�	ay��_����KjpI�J��,�+���hL �D�]�m�8r�����`]TPz�]5�Cpwu���cl�����v���ꃢ`��V%t5�0���"��E������Sd��Z�'��ϫ7 `�'zI�ɯV�<�s���G�)�PTP�z�'V=��fΗ�C��� ��7�x�uSPC��
�?I�F85�FA~;/X��W��b�%wә�HJ�t�W�<["���}���:���ׄ~Pa�%�p�S��ϐ�z2�n	T�$�u̀C�nG��2�>\��7I3��\���8E�s�����QX�D*#i%��7�OH��kp�O�~1�է#�"�p��1$�stb�Gp�ꎢ7�*;��>`���{�R���'�ʺ����l����?B�Zj�s�N�<�IT�<F҆*x1�<��ۯX7j����
�$�w��|�l��.�	�J���l%���]	�!�QR�%�4\܎��S�^p�6t�g�?��A5P��
�h�F~'L�.�èsU��H�6��dG���(���'{������XƜ�Jt��~�*���	��bJ�@��;��
;�u�>���n־頤w����h�4���"���*����{�S��1&���B�����B�)�����J/(���
�G�_(D�}[�(5ꖐ}R���_
ʣུ�ut�P�+M�{���5�ɫ�+�SXY�~р�veƲ�n3�w�
py伞�M�"Zo-PN�)�N`�����?���`�mt"����2���q!��k$��,u�<��)6E�0^-@P�e��ͪ;���NZ𽛍����i�?k�J-[D��ʌL���m�9o�e����:��S�t��/Z_��7bM��3
���ʂC6@�}���|���y���v^�L�3�s�Se�;�郂��:2#ì�`���Z�	�����8Oo�d�� aņ����]W���0���!'��~"NCuad��Ʃ�Sk�=��F����z����E f�[�~6���UY�2��>}nFS{�T�Hن�#�.��)]œ.ªP7�l�m9�G6��4	��Ҙ�סT��%f�+�a��?���p����5S�l����Ot>��7Oqw�ˁg7�ۋD��BlRP�V8�<o>��X3;�r~v��u�6ȚX�b����ﱆǯTm�[����62�		����v�M�{�˪�R���8h@��DD�Uм����~C3d��5;c��u暳ѲZk���Dg�.<���BT�WT�D�u�3��(O�	eb�2�B<���7�Hڢy�`��wǥ#��K��K�
bֹa3�I�~�篥�?�K��i�%��@9%����[�j��<��~�ES[�;��=��y�J�d�&Q�=,F�u�%`f+a8����xF�|Uqam�~���UF�	�n��4�
[9�"W����a�t���S��M��1
	q�:1�Bb8*m��X�)���Ձ��������i��T{<p,��iӜY�.����؀c|��b�\������Uz FE$����_^=L��m��6���B6'{z?K�b��/h^a�VYr�#�D~_�#��vb��R)�q�ǃVn�5����:y1��^��>9�����XD������F4Q���_kB|M:�QɎ�E��h[���n�׳��5H�e�Z�9%<��ݵ��B�9��~�g�"塰��B}.��n�@zT�JA�0�]�	NV63��M�3r��=�w�M��%�~�`I\
��ך9$# ���8X�)X���Њ�Z�^�찭>�%�7����O�����������S�h�7����a�(v^��-%��,{c�{��*.�/��^��+!��@i|v�:7��=�쒻�\3�����ǅI�D������ՠ��t���AǓd�T��2uZ��Ÿ�{�-i0
�YⰟU�����n�c�f���~5��ӗ+L�Hh�|��hX��v���(
�S��bJ��"_�Y�'W��'�����}u��U�0�F4�w�_V,rV���7�-
p@�z��!�C���9E]�N+3}a�d�Gn�B���S�p���ȧNT�C� ��V&$R˗��8#�� ��(>j�z�f�ᖞ�67<���F�9a�����Y��C�>"{;\���2
�)�Y�:F6ߥ"��<x/�vT��d��Yj~Qt�Z`�^��	��H�U������\��n�#��� "��0%�9�����Zy�����Wo��g-8�����N��S��&fQ�Ojc�u���0����q̮���.��WbJ R��!�7^���ܶ��	�y՞�w�����=��r�$�ʀ=�f����l�٥���rm�be�:vѕ|V^�RH��2bC��S�q�:0xr^Uy.=��q�=�o��t ̸��|~��N�6i����܀Y6�6��v|#٨�����va�:���^M׸���Q\l�Aٞ�Ħ�Z�Cr���U��@�QC��+��y�{Dd�:Hs�[��4�m!I���z�	 �p�S���ƤO,���qb���=�s"Va�o8�gCw��2��c���:��ؙ|q��,���.���*"���A�Ea�|ӕA�XUv����.�L.�
nd�iY�pz��W{��SM����\d�Z0�g%'� �cľ��W��Y~��,c���Z������GM{9��\Ā�˨�y��?5�Id�G�݇���j�����@�|�����j�����s��v���@Q�~Z������E��[U�{��0�J�3w��i�� >�yhd���R�D؜1.3W�6��SӷSs��?1�F��8!��8�V����_�\������aEtŒ��f��\��i�V�m��nNR2�b��+�&N2צ~�]�A��[X�3�7Y��ن��v�=a�PK	�@'/ ��BT	1��������2k�+
c{�9"�����e��8!��8�Bd��@�'xv�*�ͷusj��jn�$5xab%�x�*ˮ�n�fkh��2��ip�!�č�Z�p�����9���=;���M���Lvu�N�fkba��PI����LiL��x-��
�7�>� �y�<f\I�ò:r*>������{MN.���u����2�o��5��dv��/���L�okPv���jFċ�M��OisXF������a鉝IV$�	�y����DJ�:/c>q.��� � ��x��"	����Q|D�(D>�gї؅b��A���!1p�+`��W�;�I���j������W�7lL�����q>���Yw����7�$��)VR��(�����M����m�]���G��p�u��Z�6/*hs��_�dt�M�z�Tf@�,T�7�l�LM��.t:ѵt��v<wyj�e`.r�?K��X��V<�D����m������;�.J+��Y���
���O~���̗ �S]B���9���P�����й:Pn����� ��5!�M����k�}?�N���j\��gf�O	s(RU?,$�r�+���?:�*�,R���,b:QʛE�m�,a��ʹ[�q�X��vYQ�Ø�O����==�y[��C���_b�t�oR�Ė����=�ᝒfk뢋��:Wc�|e(C#o-U�X����dԷ�Z�!�P��ki�<��ԒLs��.�	��t�'�L����,DM�$��؁k��	Q ���L|��k�17������ t�5J?^)�SUl��S��)+5�.�YiT�W�ɱ���C�x���� )~A؇�
�R���\Z��6-���©�*�]��&40���ՖQiCһ��ax�91���>^�Q�HC
r��0:�o
�E����G]�y���ȁ�<(62���餢�w�]�`x�mj8�H}|�n%�ԎB�[��ڊ����
���L��մ:w+u����u��q��6(hh}��j#i��;��TJCg�PW=�~k ����� ��խ�N�3Hj����٧*����j+�	V���g�&fק�ɃTۤ&�OB`�dX���_���\������`"�*�ʇ��e�	$�Z�Ђ |u����Iq�F�s�I7�� ��	�Ty|��i�"/�<�,y>`��$b��\�F��K��Wf�3>#Md��'�"�q�ⴀ.;{ �
����Z���**��9��ؗ�ɻ~�		�>����Ӝ������ε2T�%_�o$t�1Nu��"JB�۲'� �KQJ1ь��1W�#߃�J�ztvݽ�̒<3�a��c K'��W�7����TBxSP�X�SL"��P�W��*
n��=_:@��b��C����s`�
dս�jww�qӖ]�Km0�\3"�R9�g��)���])n��q�A��/W`[wrv�FD6w�QeH��ݫTre�&���yH�G�����k�O��g˶���7� ï���"�֒�E�$2aN��r�����
6�[!5�;Wl�,�P`�r1v��8�oPQ=�P�S��Z��V0U�X�� �F*�3ȧed���^��t�
 ��t�H��x� �L	9y&���D�����A�r�/0�d(5��">P�'�њ;Ĭ:�C�GXk���x�������wƦ|R��/�$�F<��������0��v�B�)����	~���#��9����`�.��-X8�x�
G�>�	H�����Tޒ��W'4G��*o'c�h^!��5�?BG�/n�R�
�F�AA|#��&,��M�u�t��bSYf�d����:��C�>���>�@�e���n00��Y�$T]`�v �v�:�<��P�>���n��N7a V���h	��#!�￱��]g0+�
��ź��ͰF^��|�Z�#���l	�<�e^8ӏ���bk�gm��@i��Z.dǰu�V8�,N#�^ɦ����.��ޅ@���q]�� JK�8�g��̹�}���_aB��M����Y���|Gjm. "G�X8_>i|��y��
Foesͨ�Б�vl���E�a*@�U�~��|�$ޤ̼^#�-�t����g_S��Q]�~���X֧���ý#.��eG4'w.i�"nYh\�2��Q�ɥȶ_˻��҄���k���B���S󩝝��`�-�#�d'�M�1� ���D����οi�ev0-S�|-"���ϱ�h�;#>���r�u�	`�Ǜ�Z]d�a�'&D��5D"`�bi�)�`n��nmP��C,��O���?-9ʲ�.�}��j�~��m�� ��;D����{(�->��FJxkK�����ҏO$W���.v��&���4�J���5 %;�/��J�ʻ���AǮT�Qw� �hHFTSc��f.�/��NP��`u:}t:\N�ry�E$����w���K���O��11�μէ�(,֟E[u�������^�=�Ϩ#�6`Җ�#��<��!�I^˄�>����lr!���p�5��H����I��k�|�y����ի�&X��|��!P��}r�K�9�_�(|������PKF�6�C����=T	�q��jS!��J �����W�Ew�F�ҭ�w ��	Z�+��1�}w4+a�Ԁi.H�4i�O���(Heq5��f�g�'RĢ�����v�-�"k7����t��b%c�����$�!fv����P�>@aCa"�����%�����+Ob���Z��5wzS��X���m��l�ND�|b��ƈ��ř�FP����6�M;���*����뇼	�WA�%���� }����]���Rڥ�C9��h1�|��v��c�yX��wFJL����?�+DK&�G��'f�r;��UQQ�������%��Ԛ��d���l��e8�ye��\N-��/���|O��(�ci��R�;�N$�?�T��iR�z��׋5.�՚�'�w�k����"�=dVSs�L�6'��愺!���-b"�Ku��xSqQ, �VXkރ����-w��FN�ݮ���=CJo�F�jF�Bɖ��d�H��}�!D���[������jw�J3�[̽!�\���c��Q���4����N�u�8Ԍ�SdE�;9�P�.�]�oT��M�Dܣ�^�xA��Y��S���
�$��<x�nV�����,�P��c9�WG�N�Y�(w-.���Fv��\��Ia�a,���V�#�&�fOZ�k�_)���/�2L_�T�XX��ͽVL&A�o���P�A?�U���-M0h��>�U�(3%�Q�,��|_QR�ft�O��ڤT�d�q�pM�!�>�N�[��A��g������h���N�L�hvH���/��H�r��({�(\��5��D<�R�B��lHs	���: ]�db�bN���Y�^2X�+ �
ihy4��C*���塻��Tv'{���8I�-5Z�z6keI*7;Lߛ�b���Ϸ��Z;\	���g��ih_�L���oh�R"'{�vw���d�g�,wv-Kd���Y�:�k>'u�����9+IRL��6�������G><!QL�4l尌MO�������=�eC�V�8��S|ym12���w&2\��'ؖ}�(�U!\�eێ����c�t��w��~���4R
�[��a�#��4�L��L0d�F�aH� RᏂ�B��O嵪y����]AXPF���r�H�q�Podk�FD �E���Y�L����Px-e`)]z�l�vyо�_�W�)B�=\�H��9ZF�uK��k�_�I�? !��؉j���Ip�^-��!D���?�t�\9k�9�1`�ip��kpª������^��/d�v��/3�~Qg���pᛑK�/&�B����C�s1Y���V�S���3P�e���B�/�K�낕����@�<O���(�2��\�U~�o�{�ȞX�"��0��������&��A���cE��`ɲoEI�#A���v�T�����/��ߌj���>4�.��N���o���Ň����dyg?�!�蕑�����!`��'�ytZ���8&��'��8�(�7��|)���2-���%5 ���4��)�]�ё�n��;�������OQ3�pZ�E�~r7\��~�G^����/
��AY_8
��j���Ќr�Ԃ�k��.��DR��*�[��G��2餀L5��qh|�N�g�� �o������V�����.I�{�^,�2��c;���7MA��&�9]��:pB	tl��Һ'[y���3ۊ)+�(�p'����ys��/j�*��RKK��Wi^�^�E}g�!.���0z�M��/G�~^�0H�����$�����O�醘eSu9{�����3�uEU���+^�sN'HU$����((f���뗑��O�/@��_�72��>e�-���]ؽ|�p���U��a[�|��%C�VyO�����aO��r�H-^;��IZ}�bĥ�����;��ĥ��"An̏"�*rwc�ye�:ipK,�׬�&6o���pr4���t/���|-у���(qeJ�L8��`2��E��8"b�{��
?�	#z#!G�;�Q]Jã�j� ��P�� �}�l�5�O��f�|�N�""�NJX�v��l<��(�s�3��g
��1��9�~U�aM��fbj�®B�����x��˱�e��|��K�&L�{��nf\f���9��b̿q��`��g�R��}wck���p�Sս�(y����{�2OU���(q��WrلN���#�FP<�/�"���Ђ��Ǩ;�bΝh�n��d���}j��ε#��y��:=��?��h5�iU�r�,d`�i�*	�]�S���-�D� ��85.�� h�ӂ��܅�?[�f'�=������uH�d����7��Xu@�Xp7���B���%>�Sy{o�𩽫8r�n}�<%��)��b�f�X�٬wN�3O���YbŦ��0	zy�0@�5�ƚzy���P���`h#���^DZ��&�.�)_=޽������	3T����O�I�r��#�D����)v����Bw�C_����=��M꫚t)(�d��<D��ebA>�Ў>��i�s����ӻ{��nj�9a?��TV��|�*՘��i�����fٲ�:1�P{<�����$�b��G�`t�j�b|`�DU(Ħ Xi��ʃ1��c$n���B�@O/���q�w}���)��U7v�Q�u�c�5�+�z��%O��W� ��c��'�{��t�ר����}�R��7��T-��hOA��,���g,�~�-w��LmCk2�6)֚��Կ��P��ʱI�B�9v��"	�}���K|� 7��,-�S���b�b��^���~�[�x{LEJ8�M����=a�����+t��{��?Ț�$84[m��X7��.�7U��Fk6Ж������[D@�+|c�.Q�1��+u���O��(`���q���`��^���t=��ԍĳЂL�8D���{��'աپP��r���_���E-�*���YT�^��{�����8�@��u��'��8��]��5��C\��T�v�����;Luo�b��^e)@�[q�^���P<������lS�t~z)$��z��>q��u��=P�Q,�] �ox���r��!�$Dp�O�ܴE�V��jN���ݤ����}��Jc
��Viz�0���y��k��:��o<U~�!ׁ�+� �"������y�O�����5��|6!BUb��B��Y}�:�p��P#��Ǥ�:ZV�$rs�[�!7t��K|E���έ?>����8��-,�h0�%�<�B�,	�!̳�Ԩ���?n����L��R�����%f��t�Y�ש���\��Lin%k�^��y�$|`�$�vO��\6��y\2{D�C	�O�vHkݯ'Q�1z/!�����mD��#P��$�ޔ�C�j�	u����e��7�ߊ�u5Z���w��k�E� �6Y���"ϵ��n���%���B-�Zz	��eZ���f:��3�����\�,�p��V��0�9B�5�ʲk�MN]^���wV�������R1<z<�}c�:3>��rR�v�g��;��k��G'q�� u��-ʂ� �kϖk�i���j������#kz��$(���{>.��?�d%��bL�.m��W��A�8���W��	�����h��l�$����'dt�sj���4h;-k���"3�|�r�k��6��p�@�ћ;�ڢx�c���Ik���t���CI�F�NRϥv��f&Ӑ�&�(���r��?�Q��{��&:B�A�;��#��]�Dh���6�C.S��H86�2�6�VC_��<xC�<��(e��˶	6ˈS���J�XRf�����O������5�J�X�>6�"�k���S�Ƙ�Apҽ?p�cL=��k��U��08�M�Њ�rf�yQ��$��9���b)G�Ai�g0�l�"��_݃�O�l���t_-T���Xkr}��Ѵ
�A&�ʘ�X���˅�6G������0���#����ȓ<A�ۭ��u��:d��ڟy!ha\�1��)�s��˓Rd���&2�f���.��#�m�٬��r�41����ovC!.y�?�$�i]g�����|,nO~��H��*G"��nH|�����ꅏ:Q�y�2�=?�9���E�N�z�/r��A�|2��'I/����e���2�����_캶T��K��~�+�����(����wȠpp���|�&F:��i�?7����_^� ��}���,!� �ؽ�#H�M�w�����Jo�a8ߦk�����z�e��N������$^��
5�{�T�hȊ��6�JٸN��.�kk�K-q��~e ͸����/^	�q�����]
��6��}�y7�S�w��a�� �Ū����_�.�C*���BEpm�ooI9�m�Q=:[���I��@.�iP��F7�B�sw��LT�0 ��<ǒ���2�F�pߚrܑ�������	9�f]!^�yqn�~m�*�SW�
���r��,����XC���k	�T%NCh�LC������?�n��D��[ho۾����6���Y�%#��W�<������~+�A����2[涟����j�'��?����5��	N�Jc�ܷl�GCU��F7{ȭ�&�Q���h�� ��]b�O	�d�~�/�.���Ւjs���tU@��^�2⯃�2�f�A�:���q�z1z�Ϩ�'� ���B���|�t0�*��.�D*�k80`��[{����;9����3�C��,u��M��_�b�M��6}�9�l�2���F�1޿��ϴRC��f��l�J���&�"���	'�]�O��A�/�Q��n�R��e{�4��\.d���t��cש�}����z��~��V��}�"��=�qo����0|��[!�q(9�k�9) �7Z4l.=;w�w��������2`oMX�vh�E�.�(��7����	 a3��<q�w�[�IԀj��4:w��@?�[喵�䜎@I�5Ғ8�2_�l($�Ǆ��%hM?���.������ƛE��h#m��֣�F��L���p����3�qH��p iao|�)9$�����d�Xd���p3�O�r,�. t�ѓ��F	��q|&rϭ���RN"4�W�^/���+�>�%����ԃ��c�рS���CF�?O�w�K?KA��c�������uC��Wf��ЕcL%��FY<������-mD��n)��LSRM��[ä�[�=>�Mz*���$��|�B!,��=�P�/>�Ud���񽡟OM0���S�zY\�|�:h���쉊�¢D����R}���4���BE��Y}l��E�IA�@AR�����u�E78����μ�f��B��J>�w��Q�_�5ls���ӥ��Y�i���ICF�\�,&�Xҗ��V�F:VO������_�b�kĞ""1?|�
���r�m��\�.�:o7'b��:��(�?z��ݓw:��(�ފ�IA��w�g¦L�0z{�>�F�ݒj�m!|@�"&�sܢB����M�����V���W:���J5!�h�~�Fm1ō۽\;�%�L ���[,*���%�MuR>��8��V! B�Q������os�vJ]��a�\�	-,�cm��ʦi\Ͻ����P��RV��8�

�y��e0�u�D�m������K(�\(��ǲX���*P���o�����*����GX�PCoۀ��֋�f���;p��I�<�H:u�%by>��v�7�?W���ِ?C�}I=��kd!��A`
5�p?GkY⠭I��������e��;ؕ���K��0V�kS�
-� �g��3cw���\\k��Џ{�ڤ��t�
�ª��s�4�[��զԝ�5&}}��Fo.���}�'��c���[h�5�Z�y��W�c�Z���.N�y��cw�O���x�}��#�=��3����������gk�P&v��0�v��a9���C�Xӏk;#�|����*�2ɭ �tcՋ�,��a*�����56=�*��~�����Y����cѽ$��j�v�7�~�G�#�7��nZ��WOm$��W~̍q4z�"METQ�?��㹓�"{�4�Ա��7R�r�F��vs4ģ��2�4v`ܷ~�h*g6� ��:m�;'4��P"W-����OL%�K#��ڹ�����c���š�!����<#x��u.�N���T7>�ʋ��2��6��#�ʁ��9� opz��r�$J6n��:�h7�"��m�U��#�R��p8����9VS-���^y$k��X}� {�*כ�J��:���X���s�>^��g�m�
�q�y8yiPf�C�Kؙ�NkJ��3��)�u�V�s�^��D�IU���Ȳ!��a!Be�g�͛m�44\Y.�G�Z�kZ��&XMSES� ��OЪ}��L:܉^�/��K%�m����&��a?�?���Yb�Mqhb���&L�;y��i�{�/�q{D�Ъ%�[˧�E�=�`�{�)C%?�:���ޜG�|��nE���A��綐L��zݭ��3�O�X;fh~jf#ch^�9�s�EZ�kC��� ��x�SO�B,��s��V�[y9X�a�x��f�_$!N�,5��-j��F�A�{��W`�=vGH�1��.v�r}�x��@@b��>?�%iSs'C�`h��.?�%����a�G��q��|�!����2Q���̋q�Q$�PS�B�Y+���N��T��9i�U�x��C�݈��b�T<&K�$7oո�R[��Ԃ�����b�Q]�%H��~ǀD.��a��@�Bi���x�4rڍc����g�vi�7q��{���"B�G��+�l��D����Wч���d�f�c4�f	G��2���"0�� \�P��V|V_u0�+�a>�]a~�#t`���Ʌ���D���ɘ�Y��q6���}�"Z8���OP A���W�~3d��*Q���@�� @2O�{a�����r.��&Jٳf����G2 ��QZO
%�S�������e,�lE����WJ�Ƙx��F��?�D��U�u�����.k����lkb��K�u0����
�1?�����[?��X~ ������贃P�G���[�8�5:~�L�OD� ����j	Y���ߪ�ͧ=���)����h�v�nD^�\%�d������,�J�[����4�uJ�2ǿ�T���l�`�7�W�𷐶���ޥF���]�.��A>+�G�Ⱦ�'�@W$��is�NN-<�1rzܧf.���᭸
A�/=��n�;l����J�!���眽���.�?�y�.D�A^�ȍ4���fU2�t����Ω {�-�������FE�|"�ʚ8�6Y'l��t���)P}ԯ os��jm=�h�H�B�14롧�t���1ڇ�JY�NҀӝ��$7U7�+�Y����_K��Z��`V9� ��
��{¢8\�m��6�i�pi�-x�g�]U�#��kJ��q�oO��?+<��S���[��xO�k�mn��H��A?+5e�l-�9��_]�?��7ޫ���e��
<D%���ӟ�@�VQ�Sĳ�s�D�T�Y�Ԝ�G��ߨ{���UyC}�$��`�S��}�]��1l��4��%ߦ��S��T(���@Ħ*���c�yP+Z���1�����\�t�8�������$tv�Ц_n��g����	��71�쳁6x
��_J���킳z��iC�=�|�3��\��ϐ��9&��@�G�Tv2Xv7l/�ܿ�KݞC<���ׂ�VC��-�֒�znHC�#")���ܽ�����7�Xg�W���Q.���q�L�G��Vbw
�T����/���G�"�lc����������1�j�O�S���Rqw�bC$�8g�;�RfVp�U�>fw=`��%�-B]%%pඣ�Xa4�k�����n�V!�=�z�'s-�8H�NN1J�Z%��d���L5�Q��ލ ��6?�pY���.��@=)�d��V�^���g#Y_d#]�Ј>�b��[)"����b[�8�t�����s5y����	f{}�48>m���Z>.2��ˊù3fZx&���;8M�`;�uJ8�?2{��׫���\��! ��d9 گ%�j���<ϣvj ������|�ߛ[
��]�Y�<�����R��W�k���H�����H�i�"���*]-�����Őf�z��!��2���3��UGs��j�䱸O��z�.�Np�9-���h��ngS��{W��?s�-g����c����A	���E��D��caU���ә5�ɊqLXoH�V��7Gn���c�x�O�`�A���M���%X����T` ��ExER���OEG�dٕ]��x&��äpM��O'�k�hd�[���MPK�
�������gkJ��[r+`A�}�;sZ:C�qx�2�u�)����jm�R��Hӵo�O�ۺ�;,����M��\'������I����)~ U�0�%v���`!q|h<���S�V\U,�qt��X
s���LB�$K���kd�zp�ꟹw��B�4(^D�⢡D<Io�$�<��t��C<�$!	xڷ��g5��b�ip�U�x6�k:�pdvzq��_R��*�j-��,Ԉ�/��RX�sj gJ���vu�ºY y��Z]5���8�{Y�&J4=W�V�EGC��o��B�٤,,�]�Hv�1�UI^Ws5f�
�:�������?>�`}�q�]�h�ɹ
�ϋo�0g��!�[tu�������1��9TȀ�9�p�������D
"�h�����n��Є�*
��P�wB��3��|�~�_2�{W��|M��g�f��E2��o�1��&�3�BҹK��s���trU�q��[4�
�'Q�cCn�Kr�j6J�6h9�	��f9<A�#J���W��<��5�ݑ���f.�BV9Fh6��vzn������,̝�Sl>P�L Ĭ�݆Eͳ�~_v��WxL�"|�@M��0g��Z�Q�nf�{�)�3Ȱ�`�|E� ��l�����I�#`�*�Դ]�	�2����"�඼n�7)4���J.�6�h/��7�Sf�޺����,���
�z-E����r��w
_�V妺Gׅ���[��(��mw�^r������`�kwA K[����}3���dX��\��1՘�V�-��na�w/���ү�*>9,܏�&X�u\�m(�@"�&�:xU�i���B"q)*Q�N��)w(c�t�n�p��Av9�%E���[S�5��,M*xz�z��$v1�xھ�Q�.�ߏ7L��u�C�Ī)n�~�tNM���(�pR����o��o�aX9a��?�f�}v$9������g͏�v�ͥ��xz�q��X;z0a�F�?a�sy��vh7]��~[?:�g-��rZB�^}n5�����Fx���m�UQ�:�>���ҭ�4�l�dn��z��B��lB�%�-�t�<��x3�F\���9�޷����9�:H����F��/�
;E������r�R��us�v����Z�R@���@���!r�6 ��Gy�B%��K	Z`�lJ�b��f�������cx.'Oc0>�eJ���m �-����u?��s�0��h�gA,�~�-)�0�'|'�x�{4D�̤?"1�q#��2*)�k�[mq,���-Qe� }j��W�	;�)������e)�h�W�MK	�t��j�¥�=�~[��?�u��[������z,>��"P�It��U
��$-��\��w1W^�p�(H.����RMᓇ��׸%}S�r1�K���]e� ���P4l5H6y��yX7���)#Y��w�,$Y�[Km�_��N�o�\���/Ut�i�j�����t?0��� �D$o��E:6�5N\&7�L�Q�	#B_G��-�qq���mmWMqj����an���d
��< OT������Bt���%�Z3��o�g��z�hXs��0��*����|~�����ۢ���d&��-Yn¶��穪"p��~~�SWH�	x�����V>j�cѴ��;���H�=XvM�s���?��;d��1��;G	[�W]���Γ����M���ɕg�6��,Mʂ�urVB>fƂ��p�C �ӽ�<3���<���뻀�m��K������򁀦w�ܨ�7P��J����	�L�-d� �3Q�6X�4h�j�~+/�~	5�/�tp��K�63��W'�S�y���U{��[�74"Pc�l��"J8��oq��BMO/~���Fӳ��R�$����(�'�+������tj�*��9��HL�GLZQ���K�n��R�H���ҳ��@��0�Z�Ne�`��U�pho����0�WZF nD�`a��c�D��)�!�׫b�����g����~�\��4���fL��o��
HW�UP/��
#�<l襺��q�PJm�i�":�;�s�bw�B��z�֬�LY�.��b:����	B�m��6u���o4��������[o��P|�s>�#-����ѧ^f��2^�a��haWŌ�bx攬�$0$K�EG�o?���g�ʪ���р�����:���	�D���ՒU�v�o�䶣�K7�j;�RF�����-AX�2���C'd��$$5n�����Ť���*e�����s�bO�Tپ�hO�АG텉�I%��)��ȫWw8��n�,^UK�&#���Y�?�4�`\�)��_�-/��	m�'�JQe���0F���$���c�۽R��&�m�?LG7�}-a,��+N4>O
p�kVZ��/�� �Wx��$��O�	܂�*���aLq<9�������n3�vmO͠��^(H �|�!ݽC�#� �#��#`�>|��\>ۣ"{�A�E�7�F����V��c/�;VX��:�6�/FF`K��̋�<��ľ��EA�^��J�*��s2�����iL�q�LC��VE���"�P0F�NB��$0\�>�5�.fXa�҃j���Sm�Xj��&?z��{ĔH����t��3D�GP�n4�)�R�%�X���f}��gk7������=���
=d�^�+>�CQ�F7譮���z����D���l;��W~��=�/_Ꮓ�����^��r�T�JJL� f� �5Y���d���/�<�y�F0�E��z�����N��ZWԛEBJ������b��"��f:��Mٕ���[5��B��`0��o�T.��� ���n:i�9���*�+X6�%
�70�?��ق��{�K�Yh��4U�U�a���%��R�^��
�	�����:��C߲�ӥ��AW�S��BB�6t���̃�t�6�Gg6��FuG�"��Ee~αr�t��|�����\�����^������r�#34K��C��@w<ާ��l-rg̷\����Q�)��Wö�Z`{	�&���L9��u�ϟ�&�����#�+�]Zq�sr�Ì � �/�]ȗgF؄�PD��E�i]�?	4��\���W��I�^�7�D�����Rh'���.��h����h� ��:���q�+Rn����p��8�����P��~�s��MH�Y3V�`�������E���H���յ���j=��ۮ�a�{��(���)=�U%�&&�3�EK��.<���9U����0Q�[�3�܇P���cr0 _K����+��c޻�?���ְ<��FS�8c�wH���mK͔~L�C	�SrR(ҀV��30�8�7���Y!��/�s�n>$#t|!ے��J:��6o��U�u~�Ɵ��4��G�,�_d��\�8ҧ���gp��1�Գ������=L�m|�#�l!��Ưv�'!6�".,�¶g���-z�F�i��'/U�c�����u&�Q>��{@��F�?�����*�ZY��[����m�r/�8(���Z/��n�1	X�.�iB����a��K~ԙ�����`*��g�1���)�;��X��W��5j�t6�z�LZZ�f�ϸM]��\�h��y�9�a�z$
$�m�������+�Eypň����ꦆ�˼xG�n�D��e-�u��/࢛PҘ�����ф^"fvL'����?����rO�>��p ٗ����P,`-dW�9���<@\@f���|���>3v斫O���|�k��w�9��W��t���.�KO�?���u��͞a��	sr7�CV,rc"ɯ�J�T�'T��X�>��0x7ߙc:�Y�ew��օ,��<nuz϶	�E�q�w�rk!9Ѥ��g���*6�U�A��GX�)5"t������./��j[�^���f3@o郎�f]�@7�?a+k:lN���y��D�j]��}����C��'�y�4i������BA��A|&�p�HF��r�^h��y"�
j?HM7�ѣ��Y�	����xR�q�o�g����Rή�s}���6�mK�ET͙f��38����	�ހh-���A�aad���r���Y
�.9�/ōYT�l}u� ���i�����W�G����Rς�P�(N\��ͺ�n���u��DRw�a�qC�S���p��b��;r�������f�9��ۦ��L���p��)�?y�#%�6���]�@Ƣ�r��QC����Vu���F�\�e�t�H�7~lm����σ\.y�$�:y��^����כ\��H�Ẑ�n��n�V���M�a+gzq���Ϩ0�2���Ir�+�n������?$̬�3e��`����{![U�r�i=A�Q����yE��.8�/(�i���X�����]v��9���*1���!��>�)K�@�bk�?�:��	o�j�>���5��4b	^�M������n�`������_^�cO���b03���)��N���)3/h���[��_
���%�j�?��pl��r�z{e�!)��7Yn���!���'2uk�
N�:�@{K�`P�c�
i��L��;�V���-v�y�{�W�V��H����mxjH���Ό��;_�m�&ҫD+X�e!7F�����QT�<�,��?Ɠ�Б��>埳o�x߰H��Y�XSW�%��HhwVYм	�����d�pT��N�?��=e��C��5�&�����>h�\�[�{���E�y�0�Nx(Ht��6m�zk���c\�A�Q��<*e�p�Ш�!�� I[b�H{�-��4 �: *�����-�Z�i��A�����/F5�׶QT&�/3��* �z�gP�����]��L1�'����W�œ<"���O�ɴ�!R9sD:�yAb^�I �fz���@����"v��
D+�]��1�;���'���q'��4����D��6U���>
_6�r\QC�C�i�0ψu/ء' 2%e/�ø��%�'5[�~�

�Z}t�Z��J��2�q���8���ʙ�܁C`�p�u�����w�)c@���2���[M��DD�u�m�H�Ƽp�a4߉vG��|17� !&gcY�qUg�N���P�B1kt9u��J�ۗ�hŧ�4A����G��\�	i�L�T�\
��B��%7գ�q��a�j�3��OC��F�U��*�vi-v0|V��t��U�����}�
B9�3!����N9�r_\|�1�	�ʦ�$#��H����u@�c�EΘl��$h�a	D��~k�`$��f�`.aG����p������PԇpD��-���
���)o����B6+�5} 넷���gT�JKAG#a��W�+������[�.�� ����(�2�A�ש��T��|��y�(����v��%t��%3U��[ |ݮN�H��y��mV-ƹ膈L0U�k�>ck��:K��}s�C�����ш5���A{��jUK/��=��_n���������P
$���j炇�B����@�WN|����o�v����[���<���7��¨V2B(����o�e�A<�  :d>D[�^�z��W�j-9rx�Q��	����B���
f1�� tp>��fN�f���޿x~��r����*V*V��h�[�g��=<�8������4j~i}+�����ȋ��o��<���7dk��/�ͧmJ�I&�%o�.c���і#\�}��N9�ٯ�U�X#�N�&
y߮ǘg�r�7�ݨ2!V9.�hNjh0rx] ���K7c}%���k�?�]�6�LK�B�#�3�`���b���ҝr���ٵA�r�ڝ\��RG?��溤�ҭ߅cro]�wX�.��5��s{�[��Ұ�b�Lw�|���F,�g5�-f��{��d��"��9��5����XD�Ja麂,��G`H�g�(��l���0��@�>���
Q
ćy�#N�6�8/�cܒ�kF����`�9�)��ꋎ�خ��;�̶��F�n�H��(�f<t�@���a���,����
�9�WKtb����M��vH�a�׬%*J���z^��j���/�p��v3�H�
r��v7�IL��]�Vyk?�_\NF�x"R�Y����3�.FS�}3V�����\�I,�<Ł��`w��rg1�>"���R�C�ٟ}���� �7�[���ޑ�m�M���4�#1LH/j�3юۣ�8CT
���7N����i��-j����v�\��c�*��@�|�x6cҚ9ާ��#��f�Ŗ���_jm��N��
� �:��4�b��b�,��%'����:{���,��rR�NDJ�nA�k)���jlMx⟉�� �֑�s�1�1tL�=yR4�����������-�G��>&8�.�����-4�P\h���) {��q�ђ{�q$+*�Ҽ�Y׳=w�=*Ei��b�~��[�����v��@�e�+!>;K��ls�|� }"��ʹV8��y��A�r��ig=��n��T�M��o!���,گ��(��L��E �y��h�pG��3��3e:Ѹ<a&X6��1n�E�7����be�6_	M���ᇃ��"�PC��hmOI�k�,8	����өnr*f9s�m�
��f���'ws^;v���۫��wb2����&�E7����9��y�38��!��*�{f�-�k��f��ά5c:�mS�QM�%$5}w24���z� V8[���Cc���GĘv�+|{��5Ug�L&2�5��(����-�+��zx�@�Qk��Z2r������ /�b��l��h(��5C���d�:Y���0��LEa�LuE��L�@ �wܪ�9\�o�P��B)�n7�~�"F{z+��w�dT󭢇���-%�KP��5���*�Ru�����*X��h�6�w���<���&Y���D�.�ݏ�v��9�*�їMI�n�A`�t�(�US�����&L��3��I�I�%^�"�t��N<,����Q���Ug��A�y�#D˛��f�P��˃�/��P���t`:��^��"�t2�(z��N����^\��:��#=����c��,=�D_5��z�20>�y�,�zK�4�Lo���6	��!s)�j�[W�%~[���;���t�>+9����ˁ��zo�L:v��{s{lVgm5��!5v\�f�<ø���pR��(�9�b�4Oa�`}cc����arؕHO-���������p�98��eԩ�3|�Ծ�����c���%�. j9۰�*d]�9C+t�9�nN��?[��9��A� �*�T<�N/|�[�K�k���!|�%�73(��^l9j߱L3�Qhg��"� �rR����M�͹�_�R&9�:י��g�B�.-qB� }��w9K�P`��{SU��6���F�[.�o��'��g�h��<�*��h��eU(��h<AT������U�"�D��$^��+nX:��*��W��z�1�p�.�ZD0�d�mA��u�k��2T?I�-F�a6t�P�S>���'���l��qR�胵�� l[�س�C�
hVW-8�Z���<�R�yX3yݘ!;�v�;k�2�"�ɹ�[]:�1M��d=&.�m�A�N��?��:��jE��_�&!kBl��{^K�G�k��X�����c�b M�ܩ�J�t22z�#ag ��������5�y-���&���ux�ƻ��.Gd��2[e�[�ې�J����gzg6a犱*�߅9v�����s�L֕�t�j;u=-���$!U�]��(��I���fz��(��=a�O[��V���p�=j5�ZV� G�����r��Z9I\�/w-%��?c����0�	���Y6peS(q+|@��t��E
	�f���/gc��X\��D���w�P��Yq�:�9�d�+��.7�N<��Ԭ��2A���9��xx���,�8�Ǣq�
X��1؝��P��N�`�k~��C1G�<q8�+�^Ț�G���&No�,���#�QoW���w�	|�Ҕ��6����a�خڹ�',.���^��T_��s�H�mZƣ��+TU�wmp�6�ײ�Kf[�v�Jg3�R��_�2��@�ckČ���t���i�U���I��
͟��b�$��f�q�4��*3b�HZ-�Kh��Bsg��U��|A�/�x�L��$m�/E!>�@Ҡq1��'�,�o���J�\4&�׹�"}K�a�o��'�Q�o
�덐l
�G���A�f�P*�3O\��G��&���7ߊ�o�Z`V��K�a���9\������ˍa��.��v�}^}��}����ɑ���\��8"}_�b;2*��]l̼����e��t�m��}W��_9hv����߲�WYTll�&g�I(C�����xAJ�qj��UN�/�*c�9d�rA�9|Py1n���6O8�i�'�HM��B'�#?�NZ��#'ֈA@�.J���	���M��,�0����6|ho�o���9�e.8�
���~M`N�����V���S[���țz�5�t��N�l���6��Q���]��@$ ��R�yQP4���.s(Ey��E9����D�Y���{�p g{�M����&t���%0�ѝ�Y�t�%�m���D��%���2��5,���0���ñ��3~�1�,U��\�&G���t³	�S�G���)�?������s���_���d��ˢ��5(���3���k�fe�n�x�k�ί�)):,�zda��!��!d��޸An��=:�vYW�?�3��n��Y쭦��^]M��%��`�	�خ_%��$�V��|���C�:^�Pa�}Oޛ�y��	�HM��(��8�4���ं>������B���WD�V�"�(���B�Y���:�7�#�HN�)�d�N�_K�L�C���6�c2�%[���S��v�Wv*�x>��4S.Z
����m��M�3�rؖ��fc��jXLe��P��Pp��ݱ���KՊ�#�J�I1�a��������d�$xh,��#�=۸'�ݤ}�*�U�ϔ%>,�+egS�\��,}�=�]��(��A���qa�@�N.�-�d]�j4fjn��7�;3�=I���.�r�|�N��k��'�f�7y�%b��(����uL�,�hĜ��z��)��v��������� �f��\^U>p��p��`�.2W�$���>������Id�hn��Y~��=����9��T|��6��lu8\�Z�P5G�����TǕ��
��Q���Ov;��$�X� CV�~����}*�5���JH��2"vA��Ch�'���4�3�+[P$(��{�h}�����G�U���KB@���w鏅�O�	�^���l�jlK9�>��`�=ZQu��of��#��Ҕ
#e>���F���3<d���N�QZ�TU�a8	[L�5���������F�MV�/�y�z��Mf�`�F��%�KYs�i�hH�L.b��?�vǞWrT��l�	�4�b��}$}��v��<A�p��a�NӻM[�;Mfh�#}�u� մq���W��i��7��# ��9��8�ۗ��(�EY�y���ֲ�-h#��u6z��Y��ʾ�=I�j�s%7��XJ����*���9�F��B���T��r`�e�X�)�(((�=��t�>�c�lV��u���bAZ�HC�y�M�`#�GuK��Oy�j�E�e��bf
R>6M�M��9��B�8p턇�V��غ���0ee"S�q�z-�M��<	�i��r���v�\�������b�g���J��$�t�D�'�EWP�!��V����M��Y���y�=�4$8] �r0���.����;u b}��񳰥��$!b��eO$	D�_�ȱ]��d·��=sP� \Dp�ofI���	oj{]{z`��X��=��DIm_՜�.G�o;��Sm��(�i�5���X>��`��*�wO�U�/,Ě����/�DP�ZfL�A6h��0�s�kՀ�⹗� `ֵ�ue;��2��vQ���_A=r�g�o�7J"���C���,��ha���s��/+�@�����%�$N����X2kz67��3сӗ~̇�2B��`�g�ic���.3V�w縕+����%_��x�N穸�{��e�P�����D���vL�C8�MZX	���qmv'(Z��#Z��U�W{K��%�%��@���W�O�+��4�Ae��7>a<�/��\� ���cJ9cqwa�����0�31mn���n�^�.��s���*��d-��^�ܑ0I�sN�T�7<�i�E;�`���#�U5���Ŕ����4��8)��Y�=�3(�8"<�t���x��?��?V�o�]�_�'/����<��-� 4��8���n���`�����@LY}�������Lta�[fD�e�E3�Fg�#��7�kCiǜ����È�0Q� ��c�Z���ME���h��W�A4�Ѭ6��d�c�"0n����1�����^(F�'M�g�n��'q����]�>�Z
��;ن�oxc`ŁA�d ��:Ӓna�>q�j�����vs�4�=���hR��հ���D$Ǩ:���n}s;X��]�H�m/]�5�� ��X)�X(]���NO<qOQ	,�����rG(�Np���p4K��V-���ׂ%x
�Ը���r�I����;ķ!ٮ1(��tO�V�៸�&�g�xl/��+@g�eUr�6���nFt|�8����BI:=���>#f�;˸d$����$v�&�dF�� ӏ�plTj�����-R�%�(��y$�	����s.ܒ���]��p���z����K6X-�v�d�53���`y���ف��d�	�"i�?�g\����n�n 
Ko�z9ǰM����Q�q~�æ�gLS��C�h�؇GKY�	��"z�p��a8�e�;����:�����%�M}���..zv��M�4���}�e����b�حV�Gl.[��%%I�0�yM.����U������1ru�&��F���.pG�"kjn����nE�aH��ʃ���Mh'H�,i6�� ��e�蜕��W��x;��V׆L	�M3>�߶��v�������׎$���!:���,|Z%G~]��I���e��.f���C�$�c�H���X_���0��SMj�z��_1-�A���/}b����<H�X�<e�>*����{Oqs�7����d�����7o}�`v��(�]\����-zb��*Lr�P
�@��=�2̅�{p�6�<?�,�u�/�k,�/K��U�G��?���}q[.�W��`�f���2�+�R�С�`���S��gh��ߕ~�G>4����&rJ��Z���g����e��e6n	����%�إ	P�,{�s%AK��ދ�:�h^��t:�#]&�^��ǈ��	�>�ܰ�K9&�`9%rFW�����/ '�x�E�Q��겴�
�u��H��/����	���;)�3��0�9RG9&��3����No�EIT3�/u��1"JUH���T�TfU�p��|�l����&	%j����˗��kΫּ��:so��v�i��j}{�<W�%�A'���o7�#�F,Q������␏) ������`��؆
������m��W�舘`&1%�d�hg*�K��.fob��n4���>�AT�x����qd��fs^s ƙĽ2�Chd	�=�m"����W�w� 5}\t�p]��+B��T�@�x��N�Sj�YǊ{|��xx#���N��+�٢�q~=�I����j�ۄ��u�< ��!�&Љ/�A��ּc4���O���� i�*	nnr�!��+k��vh�	(cUh�s�� ,��a��uP��K\���Ĕ�N�!���0����:�&���(%�C�?��/�LZ�����W��!'��GselL��f�B@Rr��� ��,l_J>~M2Z��v8WV�J�X���@pL�'�!�͡L�����8L*y"�,`
Q'$=�>�Ð�xE\���0.G��ޟ��zh� ���ǆ ���/���q�F'�>��|3����F�"%��rIiT |I��������ן۫u	�	K�3�º��ۄ*�-���n	
G@��Pe'�>�K��Zy��I�"d=<0?�H4M����be5	��Eʢ�� ��,��ɕ�R�Yw"����lh������Fh
�����-O?U�������TX!ŵ�S��o��im���̸�ラY)B���4�i���4��c�|F� )~��U�#�v��"�b����c���8"_�eJG��5��#\����C�+�VA��V���� �C��#?w.���������/�kDA ik��[����%[���*v.��Άh ��;��	�vzu���D���۠�"s����H��6��;�,7y�	���{������E��O�v��t*�V�)�9�E7�|/��Ң)�ǘ�
������t����5Q.��;�b`��A���ƔoK���O��6�ضm���˒C�[	�'�9ƼD]�(/�:/�{�n*|�u7y�=�N,�����D[�B$�E��G�y�D3q}ocy\�
��hg�7� | !�_it�(�2��R\��Q
�eeP?��Gcȃ�p?IF�>����N�����nc��Jaxe_U�_������>�-n)���2�#`��#������,wzꮍ0�9�K{��M�ǿ1����<]mm�9���g�=lcSi8�S�w'��u�U^g���rC�pG�>�M�8I��l�����>������aSD-~���װD���a�r�bN@�x-�Y��V+��m��g�TM�ӣϲ�ȄO.N�ȝZ�<��If��<�,�3��C�?3��K.�N5��?�XŲ�a]��u�7u�)������'o����JK��4�*�+��{s���?ge�����;F�֥�(`	�gu�Z��&�[&��Y�ӷ�.�,s�=���-���_� >MK��O'�ęû=s�C�����]0v,X��M��Y9s6�C��d���d.����W���X���Qu�?y��[6�U�.l��c���P3�6� `(�VW\������+o>��9�d��2�<Qx/ܤ��w�Dmy�F$D4j \U�y�sA�./M�y���a���L�S�`��>�`=h2�U܄�ahD#���]Ǡ��u�0c�tr��I����fP���@�����49"�:xN�@2Eh�:�$��_4@ہ�Mk��\w�i�@�v!�?�P<��ψ]Jj��e���?�[� �gi��2
\W�ߦt5�M�ڷ�7�K'���{5˸���h�c�!Ouh�c�0}��A�Y���~)�Ҥ֯O���|�ϗ�J�<��e�:�w�-UDb�Vyn[G�B�����3���xn����o��7%k�#("�Y#��� �t傼n����X�E�n� �er�d
�lP������ ��]���ޡ��a��X���*W���dq:�SD*⟆��&=��0�Of���O:fZv��-� S�.)
��Gr��b�q��pA�V���ra������cV�-T$��)���Bc*(��׈bN?�S�硉(wʓc���x���F���a�^��8zA]ME�7����|�&{����k�u@�m������ �E۰1p��Qdm'��ޮO	�8A�z��t(5u��D��R�e�kZru�#=?�ڗL0�5XO0���V���U��ј2{�&��*#Q�ί�(�[�Cs[ƍDz7�-�GZ�w� A� �l���T�����d�wW/�蔯�60���8ͼ賗ItlNh�϶�&�b&����"��0����=����~(7�rcOP�r;��{���ޟ	$'�nr�FF�w;�B��\��3.M��p�S����,B�?nTiƻ�Q�JP�=����o���N���ii^�5�uKg��/��x�(�R��q�C;K���	1A������?hq{6E<���x�)'Ks_[Κk�T�aBgRk�ԍd/�gT�xͥ���	6�\���f|��Tgٿd5�>���� N ��Dy~ӉW5"��Z�StG��K�{Ge��p��	srZȌ!)����T8�~�Vu�G(�xb��d��>��Q'����,zi zaS���0���!���3+W�÷�o�]'��C���K�;w�O���w��(ǜ^�>��0��{Y�y�'�fE&��FT�,2��^�H�ls�SEo�p����^���"w�w]��b��F��w�Q�q��=j*���߹�MI̍&,�hU'�L��C�M�ih�		[�(N�W��G,���&��#j(��͑ʽEX���]��a�v���L�HO���M�]إ
;��ሤ���c�^�P;� _�ӓ�A.ٿ`[�I��j���y.K�C�-p^<���D�f���4<^��#�夏�r�(�	'�#ע�
���AX=QJ���'��Ǖ���29��Ҭ�d4�]%��:���䘫P�ڪ�A��J�N[)�ML2/�����9'�bs�q�?��k����V�\��/�Yp}�xI���0���/Ե�A�r���2�'�)o�,F��}��{��_G���	���s��艙PKW`��rjh��qF+~���j�1"�Q1�0LA���ؔc�+�$�r��bc���Y�{_�'�H�t�������E_�34��Ğ�0�U?��?~m?r�"�I�±�B�_R�[���L��]�l=�R�A�]uӗ�!��,�.W�+��E��fIt-ݽ���<&�G`��b��0�j'u!��9�d�z˛���1��
\����>�l��ږ��M��!�.I�� J�Í���Ƈ�*�g48�#�����,�H3$�?����J/�f<��{��C`[�\��v05
�h����OQ2KR'��)k0j���uh���Igdʭ����[��g���;�k�Y2>�F�ېUˀ�F"�%��rޡ^8�%�O�SIk��ȫ�&�O�6�����hS��l��Ѷg`�k�Y
Q6Y���Y/LQ�+_x;�3<ʑ�E6���B�sS�I�oI�,����޻8LY��|�ɕ�)��fS"�w�j�H��Ӭ�_��)~�fq�'�9>�CF��6����1&U.����;ZJ����-Dd"��c���3�Y�z���֗x���⏫�&lۅ���:] ۺ�l������o!1�Z9߫�O��5Dv
�3�	ܷ܁�=��-o��W��ef�]��ҖG=7��'<?ki�r:�/-�\I���u��灝M�~��0.!�5�r�n�_���I���]�������H�Sn*�*��H�����:Q�G�8��A�
k6�Dj��oeh�sb�Â|��X&mf�d����#�F��Z|n�iT��};Cs̚��vνMk�ă�ɑ�Q9Q�$�Rl|��������SE��d��D����#GJ�,�^�/�],X4��ǓE�G��N���	��/����/{�=�rV;�f�Z�a����NV����U�L�Ʒ�?}�g�_�8��Y{���?��0nMP���(u}���n��i���.���uF5��9zW���mFu��u٬���w�ќ'�)���g<������T�zD��~V5�x�ٰ�\i�V9kV�}�SӠ��yn�1��o�"�Ҩv5��������r#��M�υ"�%Ry�l\!�<�-=nі��u�Ow��w�4W���!6�hy��4]�O>�XݢE�K{2eBF��K#69y �b�{"7DU�,_�R��M'�@2�bh�gIľ��97v�t� �����I�������D^�R�-5u��$��tN�gÝ�%�G9Џ�䇐w��u�^��GŜ������!�j�ՠo���I�M�,�tX�MI�jbզ��ֳ���{K�n-�ѸK���,��D��	K�YI�9�Ѧ�:;�m����@�	/�R��	�4�b�$�T�TN�__yF�[�ı$-����2�XW��`-g�0H�� ��T�O(���2����Q�6�[���"�o<ۃ�f4�rm��'�_�Uc#�=� �7+I��m�c��Οt��aun����<�Ma:�����eT([����	�G�]�����٧���Ni��.��JKď�q�'
lYx���K�ʈ�ZQ���Q�i����ձ��N��$˥�@��u3ԑip�Ge@�9k��O����/^N8w�L��wr��َ�L��X�W�o��j��+��\�����FTX׮~�j{�8.�E�;9�;1L#"�n#85z�l�C��l �G������-��l�n�o�c�V��iN��}gg,#5����V�!6w�du�b8�Oo�]a��6���n5���Q��J�A`�2{@��E*T�V��z��G1[�ǣ�*x�_��L\�gؿG�ɭ!Q(�9��ɦ�Ζ��s��_5�x�g� N�+�������������aJ�n$W�Fй������w�0�����DV�7]anL������GR���1�Pl����K<D��f��S��:`
"_�շ���oX]��������¿���|�!�Ay�����g����FO��!I w�*�΅M�1���;�7��n�,%O��ƹF�E)��1��.�nz��j��9�&�AtoUa��3��PS�iOs��#*%���;�g�*ڪz㛳t�q�o�W��O��o
Y�Ё�` ��v4��,�y��m�)�j%o�~_Z�\���'�>�F�*ߢ��tk���I�s�����{r��]��������2�u�����g�q@���ۍ"������q���{��x�=�L�*t,_z,�K�,��-~n�vy�5<����MX��J��prB$��_^������]����v��~��kh�;�;vYҋ] ���������PB��b�Ցr}r�]�i�7��U^
��aJ�<f<ne5����>1�c�����1��v��2N�V�E�A�%�i	�"��9&�o����LӸ�WaH'�A�"����E�U�1�Uf4�Nt#�؎ �ry��+}��-MS�!�R��X(�B��b�K����L	�eyb��D���<��9}���[}=����b1J��6Mq4�F
EUN��쪀��d�~���a���Nx��zq��")_x��J >������}81 r�@�������_�Z�>��^��;���`�5��&�)ìG@_{F����X9G(�n����v$D]z�V�����^S�B��V����s.�<���i��a&��t�~k�;��Ջ�/�\:u=��_h�G �K#���H�v�tf�q�����d���ZU*�� $�#�����f⒅�?�1-p���s@1*]hJ-��\�{��er=�(�Ӈ���Ow���}f�|q2�0M ꚾ�G�a��ϟY��b
�7�E�s�V|O����`i���T`���>r�bA�uP��~��ӏ�s��B��Fp^�ǌK�]�����}e��L�%Qs�*��(�E�P��S���O��\w�I :Vz�'3�(��r6C�J��&��X���p(�1z�~q^���<���؏#O�>�Xa�e�_�� H�**�Ih���%����y���0�����Se��d&�X��ٶw��?��N�HrZ��Y2H���T�$������~E����'u��so�.�d��������X�yx�'�(� I ԛ;�")���7I�ʯuz�U0�ۭ3�ĥp�����Im�f�Y�(^ڷ�,��6���ZՁ�u�M��D�B~+!H)�[a���Ùi(؞
�������$tm��m?�j_�V�U��3�&���4Кށ־�/c�F�C 1�O�l;�p�Î򧘀R�h&�r�bJ���SEʝ1�����\���rl��r�����_��N��GƼ��q�mn�v;̯S�g/��ӳ�����{��FB��m����J7�]/��v�8R���	�&���.ؗ�x�DA�|y� l��F�S��
�r�:�f��/�8��[�YV�qjB�Mk��t>�"�Y��`�H�[�'7�i�,��P���\�g�P�;��dw-A*O>�$������T�CRB�$VP�����i�17L��S�:٦E�m��h޸+�ɐ+��Mp�j@Oi�4�;2C����~�q���;������RN?���,}�3�?�_r��9E�8>�h�����?3�����?��cޓ� 6�q4up�/^�8q�Q�7���::���Z@
��Q�-R�@�&��ߍ�o�����U��5o�ˊrm�v�~$6\�9T��mu9_Ӂ�Rm�԰��X{�N��=�hNM�'6z��P��u��"���ֵ�����US�;�ʐ��U$,�x}s)~�H��L*������w��d�[�R)4g��),� ��;�$길�X.��ob���Z�2����vO�-e�������]z�R4�R��$h��QnbHk���{���?�B����Z��A;�5�":�Z������'�(<��gF��m�'����[����%� Y���P�S�/t�$�T���y�|+m���_�jT��om+�q����$'H�Y�7��|���Y��!�zĆBf쨎VB�ho8�QMX��fͺ�{�q�ב)||o)$��aî=�f�X��P�Z��[�a��w�m&��4�ga:�B��g��n���Ge���N�>�E�W�qۂ~-/_�[+o�s�wI�.�+%��
�B��qYB!�h��н��4tz�$<K8�f�C�x��� �,�J�5Å\�EK�X�_�ߡ`�{9��J��*"K��:������f&ڤ�(o����	c���,���ᧈ���H�����bT ܦ.<&Y	ʨR������>J�tux��2��fW2�Y�v������"�,ʭ0��y+�k޾�ox�xP�L��2RS�e:���rt8���$6��D'�)�x;@S'��I��ytK- ��g ����j�G�Do�Hw8T���2Ip�ߢWc���l���%��rg�Ɋ&O r��Ro����]����� n�A$���6��H�0�,��ۄ�|5BR���C>#s](C���`��i^�Yzj�θ��-�܅M��l�i����=�?λm�A&<,1j� ���T
�ZR�f�W�������ni�dl��@*=S�Gw��&����'�5W�GYoB�8"`-���@O���� _r� x��"�E����i\s���Ԅӌ��:̄��y���/��t��(��]���^�'�P:.�Q7�;4�")��� ���w0Fz�y2�̵�2������-�mf㝕���%i������:�M	^�����k���3USx�!�Ux\�#5�W� ߝ';Z���
��đ��� k���_�K{m	ʹ;�=[U�+�?�O�'�Ԥ�	~Z�D�S�����w,�����*�'A΂��c*���]�0���|u���ٌ��w�zf��/��@�2K�W�Hn������Hgw�5ί�8�g\��{z��d�u���u��V��*���sq�U�5�Sk�D
���},��٭b��M�[�ȣ2i�,�9���#��ʡ�b��)^�u�6Lh9z���������j6@��g�Yy6��� �ֆ�O�Au�2ΐB1b�S�������o���<���B\����눅��t7���n�懈}Ǿ��i��T�#k��N�,��e ��Z�Y8��B<󓵻�o:x���Ś R������'ïL�����x��o�)�g���N	'��ҭDAa]��N�LI�0��{~9�%`f\|;����}[�ޘ4g���ˣ�ٝ��L6MU�\�Rm�D��l����M=N_F̉��+r�d9(#ꞣo�,���{�w�;�M����u�(>Tv���W�
���)��,v�lƊ�F� �b�����NH1�� ��n���d fYBkaO��Ӈ�(9����y:W[%)�������H"���|*W����e�����~d~ ���F^��٤p4V;��0���
t�`Ӽ���M4Xl��#��߈��C�����Ԛn��Q�a��yM�bbL���g�w"�­�ߒ6�R��v[�j��f�e�ʨ"���;]���@�I�5�]+���|�""n�}��`Ý��%���C!��$�At�6�#��)`��F�5�o&��턩��w�yy�~�VP�{ޥ_�ۀ(��;i�P�1�B�(�?!���aG4]�a�0�#@ G�۬�j��צ���,x�<{�=V�K3Ta�4���G(w2.�2�R��ퟮv2�է�~��)[�����?�cO�KY�JP�{�*�_nBg�ȥ�E��M����߅�i����7���3$��-Q�����Y�Q��qD�͡������a�یK���1��.�u.�yW$���\To0�@�q�d���?���сz�J�U��3�����V�e���_�Cp��aT��zF\�PǓ��h��m�
�j�|�O��oYӢ�'��ľ�t�'���&�1yB��`��@vdS&��n�!���_.�' U��IE��g����K�.�a̶� �V	F��/�h�@y�|E̴��r�Ť�/�z��-��D��KC�G�z��qJ�,��dk.' ���l
���f;�����v{����H�E��r	?IB�u6Q`�ǩ"q��ݶ��&���1�7A����c�T��ҩ���\i�݆fL��(iES[��۠WǗUA?��dؽ*��Cl���Zu$���zG~����q�:�@j8M#��2S�7�H�rr�!r�G�(?�b q$�2}SU����lP"�D5��Cg2;\�4n�}V�&raL����]`'��r	X���2�\O�T$+r	�(�"7�J��s�*Y�����|0�.q����y�P��Z�ED����7��r^ �i���g4
)�E�*��ڙঔ0^-Է7]<IDY1����G���0��뮽�iኌ�z]s�<$k�j��F^�B��TY�����Q�S�ģ!�����oNp�h:�G�v�L�����$�(s��hiH�ʖ�o���VW;3W���o��s������G�i%�����&�V�)�D�JAO�@.+��<O�G o��m&|�2��Ϸ�1Ec��G���u��.#y�~�Z����g��S*?*�q�V;���5?y��~ I(�'�#=��	[��&���O�ʘ�O�ō�:j�<�F(��|�\[�������ZU��i,��A�9�G�ϔ�>���g��G����V�R�X��_&a���MJq���k�&����vL�l�7��|�S�lB4�#��L�=;Z�	L��s��>Q>f���35�y��bS~o1q�o�@��T�צ.��=hh���Z����u��8#��,��
d;s��u(��խf����~���?L�"���)Dx�RRݬ�R�*p�8�� ۬����H��2r�(p#�SO��������P��r��Nu'��!:*�� �&]W��
�Ⱥ�Bu�ϔ���Ԟ��'֜`��LU0/+NU�Xq���u
�r�|�h�)d�&�B_!��V����k��D���������(0��3����v%��8��
�fg2�P�2;���DV~W�~ń�����ѝ����F�K���aT�,��[��T���p���8�����򇦐*V�[RWOA���+W:Ӟs":�k�].U��D��h�غ�M`r�IQ� 
�я`s������](
���n|�O���u3\�q<��4��F+V�����Q� ��՛��zr�#]	�6�*����:�`pc�Lw��S���1�Lv��<�� ��t���@~��-b��Yc0̞�K]3�0!
�>���c�2��=�r�f)T�e���
h���9�᥋�X�k�
S!m����SiT�6tR��l��i�PgU^�i���ga����8�$�L�i!���D�.�,�?,�18���O�#ij�t�kϵ'*�5�K��6x������k�Y
z�yg��|��Jp��jݩ��%<F_abCc�g�V6�L�U�V��0 �%��}���pW���t�}����r1�5�#W�yg�ބ٘��m�k¢|�1/��fj�[��Z>�r��iQ6�7�16�'� *�8.�{���G�"��r���>�����^�N�P�h5īZ?�_�jgY1��`��X�/Oi�o35  G�b)�C$�$�wm|o�|��vý��J��&��AG��FA��Ed�}y�h���5��`s�����+�͓+U�ц�w4����"�����"{�o���j��^��*�<<��tcU���x�C�&�='_���V�k��o�/&3�~�4����y�.G���(��ẢZ|�ʒG�6Jnj��r��u�h�ҁ,���}��
q��i���k'ł��Ӻyk}� 6"0*�Ǩx؅�M�|��I�oenV]�^�o�Kk5OM4�U����3E��WÖ�T=0a��颁x;/y���C�D^�?��_c5o��ڤ��h�h��3C���o�1���;�T�,ۄ�Ǽ�V�t�g�il�ʁ��@�~2.� �?^9�G�Nǔ�0�z�4��[v(l��z:+Vי�W[�~ͧbϻ�-��G�ur�٭��~�g�[.�"0�����4�h>�h� �	D����й��s�#�%-Iܯ�l`s�J)=T	�(#1�(XqDF��K�r
����]�7��8m�D?�q�P���}�y�
����@�s�*���t>��2hn�^��e�I�`	����"��ƩI���t�]�)�͚Ŧn�yg$��bW� 8ΧO�=����{cgN�Ȩ���}�,�LH���Fz��5�8Z�Yi�_4Ѣ<�y�ݠ�Y�΀!���!�����*�be+0ʬdf���/H�V��%��
��&DO�Kk���{����h8?�vCl��K���� L9�llN�p��h6�7i{��[0c�>��j��H��Ҽ��`fᮣz���}ib�p�dố��#��WǸ���#a=zj���X�iHֹ�%��_�A2&߯e�����'�%h����Yx�-������O2�x^~fǘ���gwjUȫ
r��r��;�pj,�ѡ�iD>L����M�b+&�u5G0^h%K��y�*��o�a�-.�7^�����@N�m��=| 
p��XZ�����3�&I�7�������j����fШ���	�r}��RLK��ޫ7�	�D�O��.���6�3!�~�����1��C˛pH��+�F"~ck�xb3M�˰�m|=��!�2�����v�"��x�r��z�Qxp+�0]��l�ȉ��45�3�90c��-f���*u���Cf'�z�����w�Y��<��s��� ;/�T��W>)����	Az</o�j��B�&`�a���u���υ"���i���5�G$)^��M��}H��P��7��NF1o*sZI��:��TYXB����J e�"� ++�ۖ�S`6�ܖv����O��bY���]��֙G��MG$��`ϦǀNK��G;������d���FdT�AP���")�u6G��@�Yʿ׸��o%=�O�����-u�U7�
WJX��`��_ᬩ$�/��c��˫�3�AF�j�"���c�g��ƹ��&�M>�yJB�p�B-&('H�U��
ѽHۯ.�j���k��a�h���0�q�Ȓ޲���}6N���c�;�?!l��~�Tv.��Ԝ:sD�Ŭ�AX�}B����SMc[a�:ˢ�������g�����j�Q�dE�l`�l�<��"� TX����ܲ&�q��оp2�v?�!%_����`�n:G��O9�� �(�/�loyD>L��|�����������S��h6�潄�F�s���Jn6_��e� 5�����z#�q�Iڶp����Z�9��kǦ
�>mv���Us�MPf�:�3ر�'���N移UbC�|��M�^	f$�W&�ݽ@��,�ف��t�i�
8��UՇ*�'�[SZ׫j��Px�9�T)���[�2EY2�8E�vdK�����6p!o˜�Dt�IV@�\�=���k�:A�{�wHh�Y����Jc�݀��b�F�&{�[.5#�M�.�C�wc��[�u�l���=I2~I�J҉�|k��T�^��[B���(������S���gqv��؜�Xm��&�p�$AA,�a��a��-F̬���)�o��q};���2�:�e.B�:�*�����yw�%*"G�x�n��#9�E�h.����3���N|���a\�y���[�P����~]��UC�"^�-t�n�R�zA���0�(��vۑ�,�ܥ����k�Q�FI�x�j+��W���&�u�H�hb:���VD���E:���Qל���ݹ�8RJ���̂�oѷ�Fܷy��w�cZi�}&�s��|�Fv� .�C"��7���%me��'^�/���{�i��-Ѥah���ww0���W����,�V�
�7q=XB#%:�@���o^��}(q�'D��D��
<��B�鋐r�#I�.��v(�y]޳=<�3�a���i����)t��pSv+�GtIsrCe�m;�B������A21���O��P����͚�~[G�ɴ�
+��8��^#���+��E�.Hň���ݽ�[�KT�x
��xV4p6���$�c�H���[n�>�^��ޣ@w,�3��@�/|bxn���篊O�0�
�&W���c.�)Y�����w6��M�i|�Y7�aD�?GW�[1���j�Dt%�!���ٲw��P?eׁ��#�>ҙ2R�4i[ܛ�����
��o��KB��=q\��G^��U���� @r�r�^g0�0QZ��;TYGޡ�[���෉��>�$��"ް1������Xç��M�4\��+�H�I�6P4�jz�aad��X��4`6��]�L sc[=5�3��b�yK?�s��Qu8����c:�M�N-��2�7��w�$SA>@X��ʎ>u�	UM?G1��P�tj�u�F}r1�+r�]��h[����h )�%K2�� �Q�p?��R���4� �>�{v�F'�Jt^x��*�T�d 	Q.�v��lP��m\ܕMK�-�8��!�;�M@�:��P�&v�isu�;���QS��ƶ��Mҝ�9�������m����Z�!�zt�;��r@��Q�C5g�� _545Q{�K��t�,���ƨ.��=�����wl̻#�)�?��-�FH��d�[����қ��T}���6��H?6�Gק�|j��C�A�xI���9���K�r�����i���֘��S�ߧYJ�����u�I�f�`M�*�j$D�����"_E�ph��t|�}9�"X�tB7�*/����.�^y-R��_�X����k=7z�̛�Ə5��3�����H�$���X��_�D���V	QH�Ɂ,�4�R��t��A�:`"�DX�9�!C�絃�wO1��I���jb'=����N������h�oӁ'U�����L���dT�<B,�h���H�Ǯ�{]�+��W�WR���>//��7?:�#�|���q� ��o���;��*����(@���b,�ݛ�9b!>�,l����-~~Q�|��:�	��Ŭ�3��0'$6.52_Ӎ4On����.����N�����p�|5�����,���1m��(p�/���L�^F�';H�F��g8����~#f&k���kJF~K?��h�I�>q�/��o��٪�a�ܽ��N�h�8��}��1f�vr��y��֌�Jc�6�fx>x�%��F6G�<��c�~�x�yS��Z��g��!Ȍ��zm�����*����v��4�ݮb
��8��Q��֌��偆��m��Їcx�$!Ѐ����z~\*�cf�-ޘt4J�˛�!�b�� ��m��^�l,l$%�L��k\#�_n[j�N�|�6����o���Hx7&]]B �i���O�Ա���J�!X㩒|TK�=���N��:z��H�%�o�R��k�Y�I��#�8$*�D��d��m�\��˅��h@r�ٲ�{c�e)�2wݝR����#9�n�c�^Z�D�9_XHo�r~.�,C�t�����<�@�Ad�~���[�3�γ�^�Ŧ�^b�j��K�/׹�f�p���ߥ�*�R	��'څ�4�|�m��W������&t�O}-�R�)�ר�D �kҸNc=�y��ML�[���@��3��Aļ?@7~)�iz5��m&���n��m�/�ƴt%\����Ї1!�E�Ṧ�y��@4��g���En�a0<�L�uߪ^�9�A�o�2��s��(޾K�TE�"ʇ�*��_�7��-��	��2T����b����i3sT�V0�P���䨱K���_�����BBV�)0�� ˱��M#�Ł�m+\���z [��=�nn��U��U����;Qy���_0�5/�X���DCA��Z�ɃWkEBV;�G47<�E���m?\ܣ�C���ϔ� Z1��-6'�t^'@����	���3 ��hg�ޡ�pȬ)TJ���0��9�n%I��,XG�݅�V��\���Ut��]?틶v�@��t�;֞3��_��z���n�6/�ˏ�)Q�c��@w./�,?�qr*2�0�/]���2��*�b����V�T`�5d�a˩\��ô�ȡ����Y��L��D ����w�yd?7v���n�±��8�1d�Ad��M��1�q)PS��V���j�\ɖw��:ሱ�e�k�<FF��Z��
�
?Do����շo3���4��"��KD�f>��O�1Z��6�M�@�e��7��i}U7�P�iL��cD4�,�Ez��7/�O3�7W�����d?����_��ȿ���O�������k�m1 �)�G�)�(.�/l�Ll�S�=�'���5��Z�6��1��y��j���5����؇Y�sB�e��/8�{'�A���L��?|��m�0�s���)���!F��A@�estԅ1�!Xg��� ����`:�c��֝���qm�Mh����m2A�b�F
�n���6��\bN�-�|��AX���1l@�Z�t��3�����Ky���0�~a:�28��˓ٿm�F!����A�8 �~4�pI%:!N���=v��1�rv����h���h3�3��źY#�,��o�=��{m�7Jt�vKH�7���lй�����7c4�\̵p�г�+3Rȼ4���N\PJ�+��Ȥ�������>���XM�q�˨]@)e+���S�sF�-�1BH�#�@B���¡��zP��
"�&��;�T��ZG�ת��X$�j�M�s+�[	x�SإbN|a��>�t����5�k��ړ�==]$�D ��UW�	��2����5�����˵���\�\��]�2�/���8X3��nDs��D��=�r&��H1���,���K{	s��O�t?��_o���p�)�R�G/#ĸ� {�/�J�p��y2��I�4L;��'���n5e�9��/<o_[�I�����H|�h��k�+J7@--��_o!m�r�f�%��m�\n��vA�ۨ���.�s�4k��}�+Pq^��`O�t6I1�)]z���U�����ͦ7�UB�Rw.�+����Cd���mjQ���rvc�\-��eGًN�f8�S���q��wB�݌����GtU�Uճ:s�~i[���#�����+�Ӗ�h�`�Z���$u%K�x�ߦ�3��y0��P��V�!�sA8��	.����Q��8��X$���1F��9"飪�p���^w�]_���w�uV�G����V�i��Q��2jm�,~,nS!�_��3�Gb��_�h�ୂk	P��q�n`5�߂���D�j���}����|��z�!�a�Q�kh	:� �L[�o���� �M3.w3�o����h,U���i#�3�O_���ӅԈ����H��Rs^7]��Ҝ:Z�q�*��F��^���`&Dh�/Z�D�s�)��$�ˤ��b9hZk�I��Y��@/��萊Y��q�*!�jJu1�_�JR�p��8$#�x"�
8�p>DI������F���
5����cF�I����o8�U���/n;\�<�ڼP�M��]0����i
��N-��:�	笋8s�+\���s��[��4G�R���(k��[1���G���%� �51�a*ˊ����{���S,>�;�5��X;��A��@�P>Q�����3��r@E�d3�NJ,w�hڀ��up��}�Y h��v�/�h9-GD���0Q�y}�V����z�3�9e���t,�߶�Ò^���:�Y�%7n�+�=;���?��sб9��.WM�8���2�Ə.W܃Z�3�uʴ:�I��`�2܌���`���=����6Ӣ^��@Њ��!�2���*[Rٳ��j��'�+	�p�ll#r�/�Fj��n�(a3�gޟ�7��wRR&;?�7��&G��������6R�NU���u��;�ҕԻ�Q����E�Z�g8Wy�w���J�I �đu����
֞I�>��|�$F`{c5s��%k�i�X)z�M�S&����
!��L������/r����ْ�5�I�K �����vU�^⺻���c�fewͼ%'KD�_�RL�#�����nKE�L/��Z���%���b��{�����Ad��!yf�P�� �p(�`�������E���2�x�cTU����nٲ`���� �D�����d��!2�A�;"�2�9*����-�T��uJ3���^���ҷ�2������.�������rɼ�يK{���$�	7풧�@���\���c��¿���A'��#�2��l�G�TT�!����^I 
,Z������s�-x�}|�+�`��<�O{������3��)�E��Qt�7�k�;Z{HN���^2�.�y��/�y-�uR�s3��w��_h�=m��[��R�H�.A�Za%�6}K��n�t�l�x����Sq�Ez���Շ��
�&\����Ӿn�)d�`�7�^K�	��ʪc4�P�s�蔻K��5J�|Hn����Y}���+�
�1���� ��s1�'����	R��;CM�F���)H���h׾OAՈ���,���+S�� ޔ��ʲ�b�L�KV,��l�ux����� ��y��젪dI��$����˖�/���Bt�"�SO	B�����֩�,�2���Fl�+��ǽ�1�t�0n�Y�)AYW�t�N-�!�}J�a((��ٽ�Yy��5G�wW�E�\���`�4�&>�;����i5���lԱ���^���<����7�9��RQ�����Iݩ=w�րT�.�<�r�Y���w)N[Z�W�L��i�W���Aj��@ѪSS�q#���la���7��ޫ��r�&����sE�8�W���nf����zV�w/Tx_pWޫ{�,*�ב5W���>+S�$�?>��������D����=�:1h��Vg�Lk*j�>������T��4
/^c�P��5���8��Ԕ��D'�Έ&�\{1ie��c��� ���I�U�1l�����T�=�!��] 	:��n�c��+��-R�'j	s���?@�nUR� �5��n8&駐m <�S��Nq�$]����7��w�t��v/Ե��\�b5��)���?��b��2N|+���9��X��xj�H'����V�4����pv��oE�^)����Ԡ���eD��R5`7��/���̾��{6Tt��R�AzzԹ�X� K�uQ�z�cN�\������x�`�!�������J	�&^%������M̲�@�>�^D�	�a��g�M�5�!_�1���6��ûTt���ѻ�]2r�8M�^]5#�}�ip5���b�օ����>;V��zMI�?�P�z�Z~J��I 3��_0OjB�[���7�e��Z�M?Y@&jY����C� ��_"�"�1���lշTNKg��1$�q�]o� N�;�	J��$�+��a�O��_�I>�)�-��R�XiSuo��s��*��ݍ��5���vQAO�4c�r�j��{�¨�M�E��+�9V3O� dꚚ��t,��Ȕ��w�ln�[���Kl�X�y/����q��eN�jʇ3#JW��$��<j ��Y*�������,�2�Z�Y!L��
��";>����#���Z���Q���@��/̪#��^U:��fc&Or�%�d~���#�se�l�{|-�k/ D{��asM����<�W���r����1��z^��
�^>��9�Ds$}>�^D2�#9��tJ����@�/z𸩡�Q_w��:����D.��֮�����u�z`���Crg�}$�G2&��\<s����;8����\��"-I����	n�ϝeYw~�1�a>/����b�0�W\q�ȸjx�p�L�/��q���j:���Ϩ=��Z�ژ��x���]�������_�B���=�y��:J���y��5�WS����,��D_l`΢�ǐ	�\��w�{t���.�<;�'�"Fɣ
�T'zt��y��XB�����:��&@����[d����_p�Z��.��v�����W�x�Lx���H���U2"]���X�L�e�
pSfK���霃0R�Y#����_�������F�[�+'U�lF��\B3����>����oV�/A�.��Rᒹ��?�?�?��ԡBS�����2Rպ�Tg^�?������Q�5{�ac:�yƞ
��b�����2܌�U!\㽟O�RL������.v�8�Zu�U���-P��lm����1+&n�1���n
�b�o�)Z�J���-��A&���R^�
�d]zy�����gP�m�"�G�N��{j�f_���8l�lZ���Ӝ���os�{�ݾ�bl�X�#d��Z'by&����Y��+��m�����Fd�>Z;��!Fs��:&�a��E��˾������ΩY�"a!>H�i������A�}]NC�YS� ��[�Q��<P1�7=���S~�H(��1�D즥�ks@Fq����t"�=K7�J�]�X~|�6��ZA�˯<��C,k����'�� Oi&�)��W/xҨ`���J�Um�B��n-���\4�bH�>�<��6��U`�Y{&�f�V�^q	P=�(������C۶e��pI_#������$�HiF�ٍ��6e�nM�e��`Ֆ��r�ň�����
���2�5�X������*���3����z�s/oߞ��Q�}/0��6�z]"�6��"T<�3@����Ǫ��)�l���M 8ah��G��Ֆ%{�\U?�uEL*K�q0@��5-���SKo'����'<�E��|)�VwUv8�A�&�����q�l���2��C��h�J���]��,z�	�˗Y��ٮ��51�S�
�}�T���D����mF����Kq �I�mWL�S��͹�,)�>�aW��@N�CM�`�@2��x���y���� \�����ݡH��+m^�N%i�3L:�m*Z���?,DX$�"�%�Z�B8c�`���$|z�wP���n���S_�r�d�R��������Ѳ�#�.�4��#A�d��@��:_O�P��)\�G�@7)�]3X*brM��n�f0����â`*:|�v;�Bq���ٯRo�X�ּ���.���x��7m�վ�c/�B������H����� {�m�z{Ć{D�1Ӣ/ٰ6D+�cv��֖L�Jz�#Q��ρv�h"n`�,WO5�:X���ԑ0�����jY���o���ר������H\�ߴ�U���#�LU�����m�>Q��+!*��Y���asJ���obѰ$�#H��<��n�@�[�٨\�"�ܚm�L��5wSJ�3wJ��~j��!��Qk��-pp*X�FX���๲���`/^�yOO��)���������]r��}+m�Ԙ�7��OԦ�j�M麷ݺr�Y�D.����j��j�ދ䳪<�j!�����j����{�Rr��|����,Sh��v�_c�hd�7����fe��9�B+ɏ[SNqLg�xs����N��ӷWD@T̻)4�v3Gn��]t��>7�C	X.el$����YjD���c���2�1`�jE�k�ͺ��G�F�:���-P���f6����F/I��ۍ��稊Έ�S1Pc?#Y�p�$a�F��Ȕz�� ��/7!��s"���[V��U�N�i�s,�u�n��D��u�%�#�^_���b8�F��/z0͝}crh�A�9�����ݕäkAQL�o�H�E�\jJ��Hh�r��$�^7 �2��6��wDj��0R5��=��^:��t��Wɽ�)�k��'����O��L�oLv}��Xz�
��t��?l���\]������� �i6ep��Wpߛ.����Ǵ��&xm�x�^�9���5tdK���d-��\m"�_��Lvߌ��?�������~��ޝ����\�.۸&3?�6r�.�z�s.������r�B��^��&	�'%��d�>����4��0�[n~)�H^q��ً�q�|�"m$ފSK4n}�ً�/+`ΝN& �1]>� �z���B8��cH�i�=��C�(��6�;gW8l��� ���E�R{Xz�u�-3w#�ș�1t'������� �}�j�,*�/��D�I��������iPK���� �^���p��xék"
���+��n�
��@��-�ވ+2q�19S�dc�3J�CK����I�o�Ҥm���C��=�.+���9�b��C�n�թ��آ���_s�
S�
>��9,��)~��|p��ElVKu�)&���3\N���zx�3�?d�ȕk467�A��J}���c����;�ЯL����M$&������9ut�WK����*�q�b�2�	P^�ʳ�QP�Kt<Wj�f���a�zG�� 2��#&� > $�&�ʩ$�Y�����;Ap�B٪�{��7�;g���qʲ 3��rײ�z�6��+�_��W�V
R��i���.�҄G���=^�פGyL��FF�}�<�d�O&wL�ԩ3i�Y.�m"}B`w��TS��uSK��dL����<t3dyoi'9>>�Ѐ]X�)yb�ӫ�y���	�!z�u^L�v�c�+`������_�?�;6�W��)A{q0^��M@��vK�?"�\(����2�~)P��ʨ$K�C
5������[��g�C����_��"(�7�~#Lu$!��2D'��@��l�pKt�X�h؍@a�Ϳezo�&��m���,w�+ZM"����?���%�����ξ�?K�I�w�0֣6�w�,�*�l/�^�@���*�բ"�`WQl_�����v@���w�Z����_�Q�������I� �׸�;.�ٙ=#�~��:�cp�!��\�/�����Úd�s�Y���x�&�+���Ve�> �m{q++c�:��]J()2���c������ԯ��}�Pr1Q]B�:�4/�d������	��;넷�S�u���[�~�����/L��h>J�{-��T�8%��|�!I���Y���m1�����A~��أ�����(��l��_�o��0��m��%�'1���]�bm_�A��O�F'�E��}ɲ%���
`;%qF2V�/���9����n9���?ksl���_�DK�t#O��a$	�� 3�KwinԲ$ �[]t�P�E�����O�;D�bk���@�{��4��d�s��F%Ժ\�?'�.Xgo�iD7}�����y:4�^Dyb9�itdk�c5xo�x��V�k����:鵛L0V �q4ُ��X���Q���'�70&�@��V�|⻧(E޽8#q���%��)��>�4�g۫�A�d����l}Q�hbx��b���׻*��77���^OZ�?<�-C��w�k��D��sgMD20�Ύ�mw��2*�b/!n��a�1�	�A���Se"-.���W�����@iu� �ow��j4��?:��߃KbO�H�l��M�)8�ot��m������iA
2�W�C�N����?���\�د@y]����y$�@pb?��P�Գ.�,A��L,ih��a� �Z�ƹI�g&���6�_�MR���̈"���gfD�"���F9��� ��J������ƻ�/��c����p��>`��T�8���fC���H���9�a��B�� �������Q��쎑���W���p�]O��F̡ Q�TM#�n�S��36���[�9�KT����c�������	I
�h�Ǆ$ki(���9�TtY&je1}G9}� ��z� ���/��j�����
d;3�d�վ�5���7��#AW\���� q�������jE59��#��A[�0���xs>k����
��1K����p�����4 ؊/R^)�)�Η��W��N�`)�嶜�p�"}�56C0j/T�����2�s�p0��!�ei��k���~�NV�S�^��{�"�k��C~s���7i���F��3k	�J�]�����!��*k�����VN�@�A���3]9Ӹ�Gz��c3 $-�/{���6�"�� �Y�L "j_⹗0`-�u�MW���7��A�~V
�~P��V��jIX�qͷ���l�*�`7&��-�F�\��lc_��*���S�v�.q`�O����"v8gkk*�G������d��>kN@$>�I_"�<��G��Lb �F_ќ֐���:-���O~��l�%���6x�\3l�ٗ���[��֢tԖ[ߒ\�v�WD~?c_��m(�*�K
���G�zH>�ktzU�{�g'�	���ͅ��E�� 0�Y3�2L���u?°"V|<�Af�+Plz�~Ci�S~��iR`��sƺ�z��6�Ů�]|�����_���<!�m %���
3i�5\�Q�Eҙ��8k��x ×��;�1����
S���'�B�����8��S���ݞpݝ��(�-q��F��S� �{�H��M�0Z� �O�]:-u�NoN�����8L/5�bL���2~i�h�+���~1{cgw~� �t���xr��;�}����^�+�fU#��������A�@Cb'm/%�*)L���+��,�N��ѱ5�I뾕��摶�M�����$�����<	n��G�����ب�LY����D��d8�v6��E�����G��^M▢
4���b�ن3��w�;9�n��;�r5~(���׿w�%�2�>X0�u.�٢�Y�e�Ty|(��"x#]���G"2z��p����0@k����
Ŀ'�y��3n�N߫�Bf)�i�D
��S[E)�\Q���"׺�W���< ��Uq�v-Xl�50b�1p��9��U͋Y��bKN�����1} �Z�e���D�2���7s>�WO�y��5X1d��'���i��O)�^���,�{��e��|��5pmZ����	}�5�^�-)�H��mm ���!�.O'�.�-Q�EG��H�uR��Ӊ���a�`�aSm ��K�[���<������q5��د����E��3�'+�n�[>�o���Y��6�ݭk}��Rkie� ���#X�ϩ�g����H�Kn��A���j-����E!er�WA�27E'�p$��e��̚3�A��mcN�ј�3Sm�%ɛ��s(�h�*�(��*��:B��z�=�H��ot��$�ʕ��&|'����ȄQ⋼���7 ܓ��%�*<?�|��LT���k�3��:^�/b�K�� ܅v	��6������F�T����;Q��Va2�W^..I�?�]���6�4�.s���+�� !\wJ9��f�ys]D-�X���L`��hXݳ�$OP�h��=�޻^�'&	'D�>�fn���^ݒ9:z�ׇ���	jWx*?���n�;<y�7kA1���<�^k�r�f��|h4ј�Q؎�`���	��J��x�q���"?�C�{���I�^���m���g
_hI�d9�o,0{�����P��,X>?��B�M�3_�8��Y#uDݠ��	���nI��rճn�B��?&�^u��.��Fĭ4��aA�w�%0e�V��U���V/5��h=Z��3t#�/Y݄������Vyo��N�L����`F��~BrU�5~�,�wH�;�6%>조���
�x��F�+S������#��P�u_���^��ƼdL0d�i��ײ�zƣ�������>_��N�MtX�ก�>F��<1Y�3���Iw���]�ɓE�N.F|z+����@��L ��F��L�R�j�������� ��I!xq߂\��,�~Ϫʹ�?R�'�+@1���Z�'/;��|��@��i��+���f�q&1d���uU]��Bb�s">�(|����?`�*�g�	���S78P��BE��F�7�ĝm�*���T@<���O��Ύtܑ����z��E��<�":m�O��S1&�|Ժ	������pde���a�:n���ˉ�ʛV �����s�<�*�c�tj��N��W7���2�_?a�rq��c�o
C����
	u@�Y鰔?��=y�Q���ר�Ta��R���[����l�b�!Q���T���N W�\�d�C������żS�(�gGj�GU=eNޣ
��&C:߻�]�KCΙ�1P��\�PQ�,�ύ���-�S�(���8��h�Y��l�6��r�Xl8��G�x�( �&�7�^�K��7ze��8���\+�����/>��������yQ|KL8�o:�C^E��Sz�e��~7��±/�i�:s���V9����h�j���yf�gT{�XVhi���)�K�5k����¸�����k�����|�lb���`
��,��l��j(�2�(��}:o&Ĵ��	��^m���@�mC�RLG��~}����C"�����e���;�zOE�e���H��(�嬭�<��TwFG��h��M��p�=`$h�@��@|˕79���z�G�B�1���n��X��u]�0-E�I��0�U���>-�?�P��W�zpB��{8�؝�j �FK3���.�ew"�}Zf�oa���~�q� �oq�	�z�$�?XGdrr�]�V�U*�����z�
2�[;���O9��b���Y�n�����߰aYd,��N�����CTa����jsd!�^���<��w�[��6o�&>���Ln���^t��V��PW��*�p�PJ}�ܾ8�CZj&�F��e@0ӯ8�,�f��1��G_y�E��$� ?9O�)���AwU"����p� Dv �K��7XS`�Y��5���CD+�c2����u�zĶgR�����Ŀry&���H�����̏�r��B�JtLΛf��ꂔ�^���R�z��8��դ����e���p.���И�B ��D��2�� ���$T��Qn���0Z���}2`��J,����#��o�Yҍ}���^��5>Kn,���.����K�jg`2'�~�4��L�D=��ú�Q��߶E �KnӺe^�:�#���=;��7	���� $�$A�h�S�=w�*|+`$-��S1[��{�//�q��m,�k ^�FT{���<O��/ڂ�-K/�l;���9P�d%��L	�����9Y��s�6-"�x��Gݳ}�� �д%��u�BA�/#�`$do�b%{+���m�
m�� ��:1;����ˎ�C�U�4�a������������"~��ȕH�E��k��nZ���8�-�ys��������VJfQ����:(n�D�P�N���C��Ā��7C�
M�O�Ü_�Ȝ�QF��h���ṝ����$vI*����r�_T�@�� #,�#�;���@����u<��4B�k� ŉP(}��n��M��� ���Q�0��k����P�jLUl��~x�@!��f)��l�{j�:���|���W�dBY��\���im)]|�3�L	�0%hd��bql�8��9�HI=#>��w�����5���Xom�$Qs/�՞~����kְsLa̱w�d1��8��A�p�$�3�f�i��/5`�4Ik"�V��䃆�B�g��ۛ�P�ʲ�]=��v�G5C�ә�m����M�d�=T��te?]7�Q�|�e�8�Wn�X->o!��k���4bM�z�a4y�X�ଯ� �Ohi�x^}F8���Ȳb���Ĺwi�W���.}�z9�R��kT�x&���J���o;[�����nE���
@|�#���ՠۻ��͉��F:1���T�ih#
�t��pc�hV�>J���yO�%?�~܄�gi��&�[��J�5~b �%�|?$�v�2��|���A�B�>/�!�_EH�B�l~�ӫ�6r�S��ה��d��/.Q�j��%�<��hƵ��ijb���3�v���2�X��dT�E�~�8�\g^# fD,K�َ0��;ޮ=c!�r�C`XcE5�ɏ��p+p�u�n �1�
� �������B��	ݬ>�
2EQar��d�����޷��O.��n� @l�1�����E=��Ż>�`B^{�W�|�v��K\��i�����
?�c�D>Y��]�\����_�z=���ꟙ���œ��&��E��rk�Cʶc	�����6RaWo~�E"��U�e@m�\��Ip���1���~!��#JG��7��L:'^�� �NQֳ�,s�14D�@m��P�����\۳mPO���a��o�����19
J��e����j�UDe~*y�#Y��`%j���[�����zyX�c]����"�����d�.�RM*l�t=H��C�NC�
G����B�9��6X��"��WZ����B��û�0�嶬9Oƕ�㩜J�:��q%, ����1o�ŭp�=9����:����wK��PuW�)�z	���!�3B��i�N�2��P�Ɯ����C�F�qJ�C���*�C���&�����A*��t��$� hC	��"?yMk�Pjģ$R�y}�-3�$�.YJ@��L\P4�-��$�+�i�/�1[�u��m��W��^�O����ȼ��� ,Q������?�d�D�I�"ٻ�*<�TV��s,�+?�+:߅8��S+5��cG�{�����l֏"P�(��L̽��55g^X��8�BRx�z�c�!�)�f��}�x�gE��9��n���>�ۀ��.S*.>�����z-#~��C �Ub&�!�}j"q��M��6Ҷru���(3�8���e(qQ?^ �o3;Zo��# w�gh$�$@�k�t���xF�ϛD��w�q���"�i�����r���P��!�4�+��'�b��܁�f����j$�A¿�9�N�θrf2y�9�ue֪{l�ڡ������v߯.^��.[���FmQ�4."�iX�-�j>~�%ښ7�:��X���bǹ��#�ؼq��K񥯆���?V!��p��VQM�@b����|L��D��Q�"\E@�k,��M�����鴄Ez�9��b��`�U����[������7��3Bc2\\߸_i
[�6<W�1g`%� ����6��M2P9�%��j�K������ȩd*��1��H5����7��ӗ|+�ʷEu	��������
��+#ߢ
c��&�%�V���ix�1�ô�,�#v�	0%�,)"�2c�YU�GM�Җ�S�vB &�<�Z�%����l��?��?}?~(Yp<�#zͨ����j�\	b���ʸ7GIi��޲8��Gj���V��Ϝ
C|}���}ց;-MI�Udh����lE��b���ԍ��EO��u_�cK(�{,�C�Z�]�v7��x3+��0s9�|_����J^�-XC�"?��,ގ��;V=�0964�� ��!z���2� �X7"&?��֦r�&Ol7�_�)ˏ�ss]�ե�>\єmY������Isx���ԕ��O�jo����e�ل*��(A�&������~�5�QF�� ��򗠢	 �A��&�S��钃�f;�&����=�,9��5�h��3�ڐq�&aG��o�w����ITm?�E���ځ��H�e6�f�b�1�xMtQ�*Z��5G���h}��x�V��A���w����4b�Xc��+ Dw�̮�}��L�]����A�W���b�'�Ȉ<s.����:��˽:�)IN���,�@�-L�P装�>���,�'U��Ù��+�?*q$L� >�$5���
P!FC� !}[)�u=mV��9���)�RzߨH~֣` +a��K��#L�EA�J�8iꮥ!��Y ͽ���j�!���-���X|��c�[W�
nۯ`����R[���~�>�s��}v���oS�5�p-��C[
��cL(:����ġ ���u�S�v�핃��ƀz�4Ν�jw!�R>�H��ѹ�2>�~��xR��A�(��q������a+��3Y\s�����щ^Dُ>��Ť"I�"Y��m\�>�������{ĈC]ý5X�O��6�����"��ퟀ�[k�B��0��qT�/� ��X?���ԉoa$>�������~S��U�rl�k�__#9�(�qOo�@n��|ga\5�.��,��2�Nው����!7.��:�6�*b����6XՐ�7�|�+<p-�㆒��[���:j[E�ц(��#���^��`� N	LG9���hR{S<��3	�L �`����<?Wtg/��$n�]C������X�>6�F<G����迖/{`��9+^ԓl����N֚�춖aI9[�i?P�V3F͎�`<�g-ھ���h'�p3*��ߖo��OC ����o�����ml���_���!����*���6�*�S'7��w��fp�4-j#fĜ}���G��Y���"�㣾�rNPm7is������.p�EՀ�����y�k��pC�\����P(��ޙ���S���6��+��\)���:si���-�OC���$�yw :���[�i�+�T@1���^lo�IH6��t��Ce���*8�R��8U����� �����OG�7V�z���8|oHP������Q^6p"����0.K�!�za~�a�?x~5w�Q��C�
��Q$IX��z�����u}W2�Ol0c��8�Ki��c���N��q��^��E�����:�&*�,jF�߮%�JR�~��A4��#=�mNd�D�j�@�փ F�u�p��Yw�@4�@+Z�KF��*Q����O*f�=ާm���' �
 +���:�<��_< L@i�f<�OK�4L�&��0��B��E
�2��:M�hۢ"d�cQ�{Wu��:�D��/��>���Nj����&ս�~��&������N�|m�?��3 G@1/��z�� �����a��,r4�p�u�WFy*�_`�h�e
U�Ω�42��.��l_%�A@Ѽs���R�Jʹ;���:�B������ǨT�K�X5�:�G�.(�40��	'��&A�7�0��~ؚ�]"��7�酣upw{�i�-emN�a���+c�'k�%�П�	�g_s����%����oK���+�ࡴ��ON��p!*&=�d�[����6�v�Y�6�{������*�վ�w��>�\��Yxs����W����������!m۵n�l">N�v�'Cv��p��)N��Y��!�sÐmh+G:K�n��#�fP=��7��/� ���ژ��qzq�h��NOY�̐�_Eg8�?�i�=�Wb�F�� "�M�&SMB��4��@?r+�:�j�&
�?��� GD/\T]����W��E������Ib?�E��T`�Ϛ+a���&�q��;zĢkA<�ӧ��f��Ji�M���u<������.����n��+P鬻v�63�=�]6_i�ǈ#dn��UO�m����Z�ؽ�F^)���{~�N,1&/����)�̉��)S�(s�}Р�3Z#��'6ϰW!�]��q?Z���n�.O�\ږ]�5��&Y�5��ZGLuv������l�s~ڔI�Z��)Kz�ճ?���]�&��>�2�����?N	p��켍<�t�\����#�{E�w(�!�D¢��z�JH�h��~���d����`�(`�ݎ�5$��������B15�������Xb�����m{_��ۨuN� �q42=� Z��L�Z�\/�G���c%g��n�jp(A���]�	q�m�+i��.;��!�;��~:�l�6ˊQZWo+���|6/��?�9L[�
�0]Ԥh�x#���	d��W���́�h ��V@��b�?U7��y
JB
X��J������r�X�
�����C�Y>0�B�Q������7���������'���턡�+�=�i��|�ܰ�2�w��ԈB���w���9kI�h@�F�`9�]m��Y?��[!�{�Y$�.��F�����%;�t�$�q� @:	l��
|]o�o��w\��D�%�!�����A�����6>Sn�zv�͝�E��%y#Y�������1���ƭ�Z�����t�mi���(�,��D���/e~�r�:� �� o>����q1��8�8 5�w���*y%&�O�˅�������.6�����5��KG����eD���<_��.�8�P��h>(��X]�>�C��A�?�!�L��W�u��/>@�Iwd�؟�i��;\ȼ�B�N�ߘ��l�{I��r��3HC���?p�������p'0�#I?�}�Z��b��
rY�,]~�Y�/����wЇլA�����#p���^a�Hֺ<�9���]��IX+��?v��K���3�fc���2�r?��\��}���~��5�J�”_k�"s?aO�Ss����E���x;��ü�C4��eN��{�@���q��'7�P M'}S�+���6�zunw�;ϖD�o���S�?�5��.���y��t,��]Z],*��	�m�!�y����BDX�����~��ه�Za����m]rMĊ��i�4��ғ_1&� �����B^�"�K��Ru��G�Ǯ�b�_�y�N_��.~< 4��r�jJ�J�J�'�ƞ��'n�@!�Ĩ��T=�x�Lm���к���t�����o�;J�<��hko�x$p�t�!V����o��G,q	*��/�'��?jz�������w��iȼ���G�j�.Z45��!��网
��o���۴�&��в��o��V,n�>O�e$,�!!h���	�V�\�U�ɠr*���R�^V���s,(�l%|�}S$�[�[��ͣ�U?ʶ>=R	VY{�=&|����;Nr#��h)�(ߟJ��+"%܈Xl�o(3�����vX�Y��� �_�	���+(�Y�Ɗ�uFU�N��ѥ&�.SivP����5��a�La��#�w,֩[k�ٿ(�����lxp@F;�u�ĸh�ɏ���e-f��a'맃�b8�t���� �����=����EW�q��R�s8|Km-�8�~@��+�#���T߹yH��/�M�v>��t{��J��H�s���U���'>��� s�@7b��ƭ�)Ʋ`�u�jq����X0�����N=z\JCh�0!�?4��P:ڣ��:Ԭm�T���%������ ��[s�����C}��	ɻ�P4P�m%�s�YӴJà;�&�U�� ��:�����hl��Fi|�D;�/�bp{�6ud.)g���'��V�:�&)&=��Q��'�:��H];0ca%�{�څ<=7���ӇÖ�cE���-�&t\i4	�h���R���a����";�4�u��UA_�q�x�}��E�m�Igx�nxܹ*<�<�ݚ���\;I AM�L�H����Q
±��r���r�f�a� }���G�Y�^�IS�,��]��"�s#�۪�eњ�芼7F|�dt���ua6W�͗��A}�C`c��R����Nq��
W{��`H=ھ���<��#��xc�(�
�,r����䄴�,�ᐟ����ۦ-�:��^6b���V��(����� ���D�+�At�p�74&�W?@I�P̋썿����
��S��*��"�'O`�]t�9D:�W�(_�g]��K�`
��5`ܿ�!W�m.���0���ID�^"����m����]򾮹���q��Ou�9*��%(53N�@����*��,/�V9�^� Ǭo����#�֙��wf}L��s���c���<�;����r�g�w,y�U�.�jb�_�9����p���,��	Ȕ��0$�b`�I���f<��������2�_3WX�]����DÅE�ˢ&M&y��%ժqp(�Ĉe^x��e�-;'s�`r´����H��ҡ��Ӟ�BBN{�&�U��:"�m\&n̍����l�����/�x�z��&�]�]��@��x��<���e��(P���Ja�O�K�.(b$9+��I��Tg��%��2q����|p�IcD���x^6\z�_Կ�ۨ�ȞPEYi��fp��!(TE.��bu-���#�5n����j�_���-iܱdߍJ@��08s1�d���OZ95b�`����"<��dw.�}Y\כ�O�ō��]��/g���{+�I �?ݧ�](��T=j�h�j>��djh�����|�9���7=�a�\y�EZP�o��	� 6Y��n�-*rPu!��*����7PUM�����Lx�b;�Qy���\�x[p=c(�[�N]�����Ȗ�)_z�Eޥ�8�_���&_�ӰjC"��6�*�M|�8��z�_yF����*���d�,�R�О��Dn3�,�!S'���=�)�<���B�����+�F"�|:�gx����L�׻鉹��LO�R���|����p�,�bŝ|�|D!��=�o+��FT> �}?ۘ����Ȧ�A����.��x�<"�<�y�pbeX|��	߾�9X`��3��L�e�j6)b��z<�xX!��c�;EИ�B^;^�J�k]�[��ݐn�iZ�;܄�+��J�Ӈ��U;e[��
>HY�X�`R"��6��|*o��`k������_��$R�Go��1�HN��p��
oqag����%0M@��8��=b=\�o����b�[wS�G�u���w֟^$ɻnP�o-�L�� ��.�M%�0�q-��d�(�«^t��Z;�p������۩b���2�-�Ҏ���0��`8�D[��o�+�w����*o!��L'=���tޚ�_򋙌W�����"��b�GV�]��U���;j�W_��Զ���+������*�gS�����s�K�=���FTj"c|�ٮhhl�Τ�R�e24�u���xR��s�栩 �̐��L���y��}��w�X�S���9�)�/�`��p;�?:6�DM�{e��+�������x���Y{_���ĵ�DÞ�F�ejR(Cp�x�����(^OR��^)��)b�*����'p/7���w�"S�rH90�ֈ�oM�^n�����p�	����,D1r��BM+ �ɸ�^�I?����g���ڧ� ����t�"ra�Z+��j�g��D�l�~֧�x��򢳊�|�NWܛ������yڼ�/���������y�?�p�~Dǚ�V}w�:�.�v��=ɇ�v�f�^�@Az���U�� ��g��]·χ=�i���� ��dȨg��	�Tuò&@8	��q�%�{��H��f�]�~���O�D\�É?�"�*�<l~f�d<���}�s�[֭J�H'�p�+�֣{`t������^T,z�
oOd~c�Fl�����
���Ȭ��M�(c���PE=TI�Л�bڻOw��9`�:��gɃ#W�TG^����<�V�3��D����x9	~�4s׿�؂�=��H�K|_Ю2o����U4�K������m���0"�2�y �f��z�Ԯ��+�١�woȢ����������F��։��$�3Չ��3!�^jfynz%�;�N@lGe='t׿�0:�gxb���BJ2g�q���v�N���6��A�u��?�\���Q���x97Q�0�?iB{\�����6)�6	f�{V�[]ΝB�oуw諬�\n���@t��3Z6_X]SA�I2'Ŀ��s��G�T��" ˃E&x�.F@񜽴�6�R��5�#�՘�Fтx4oR\�bz$�X�j3�
���5Evn��	�MB���̗5Y�����NŃ"��xcd�خ��j�RJ��6��O�x%�ݪ#�m��z3`E%
��Lp�����xN��Y�v��~k?���Q��5HA�":������ea�.�,���9��m��;z�U�v߀`�u��^�f�nBۃ`�f���dU���|+��X�m�7���^ի��׎�0A`K�\�q �:�"%�@}���*�sγ� �m��-��\�Mh�n�`����*�Uh�+��#B�}%V;��hwNN՘�f�
�����71p�/���ô�G��d8E;���`�el��8X���,X��Sq0�9_��|��T��Z�����Y�VX�����)��:��[,tټ_
�Y��o�i^��$+�eK�9 ,�܇�Q�K�C��=�%��Wl��/��/�+:Ct���ݢsm�bE���u$�>�<�7�ߵ����*�1��E��N�S�������
��*1It��cc��R|���-+�h�	/UeR�$4ˬ�nd�-�����K�*�xv4��]�7q��̾q���jcr$f�#%��[���=6�<q�p����0 ��h��4�e�W"T7ؐ�����?�8S�a?�2f��X�ab�.�9�!\����䮘?hM�����=/MĊ�o�Ǡ����{z��,E�}|�qq(˧�[��_Sa���Y��2����Z*5��J��?���	�H��eӯX�pzҩ���+N�0|�$���[��о�G�+�D���(�¨Q��x��,
e�#�Yc���������7��=�Ȍ�IQU
�o�6<���!/�n֪ Ȏ&?l�O
yp(HzJ:�	�K{��c m79�9�O�*�h��Z��
=���0���P�2*=���2Pw���/�S���L�y��@Jr��A�D!���ğ�~���	 S��M��!bv�P(�>P��?�$!B�O:��v~I�l��~Uu�GvX^8T2�R�|�m�/�oΞ�:��-�B�by���k�{}��Q�� &���6����@*�6���>z�ĝL�G�de���\�T��<�����V�; %��o�q��h����̨[}%�w�[���(�
DO����E�0�%��7�;��w�� ��ӭ��7�,ED���"�O-�C.�?c)=K��B��|���[��f�=�m5&D�C 9* T�1Ҁ��A��OX�˙��+I!K��ʮyC*EMѳ3���s��H�m�:�����K�LIB�ݣ�N��U�������T�OI�9��4��t���yS@���y;ۃ���Թ��bG�>W�IR��^�ҡW��#o%�z
�آ���R���pw�C���(N��ژ'�_JG샠�mt=��R����W��]�)>2�|&�� c��|��&�:.f�#r�`W��7��D_e7�&�>�r|�r���ބ�B�ɣ�A�⮌��h�g� ߣd8���T�Ӵ����u��u��� 6J}�s�
�Ke9� &��.�o���d����[�,޽�@�9��Ԧf�Ү�F���áǌR�_D�?���u����R���� ����T����>��TD
:ʲٙ�U�$2������d�����{�ԼN�)"����OKA��z�j|�V�VĖ���A�UO㮗�o�3����Fi��W*Z���M�h��C�����=��y(G���j�P�Z������z�a��"�*�:,V�k;/�4˂���b�Aj��Z�	������S�s�Nuu�t�a�A�$���6��ڻ��2ޫ�ӳCQ}���w?���V���Ԯ�������������c���'�.��#ky2��R`ټ�wI|�_��vkq��f�3Êi�BH.^^v.��`W֐v	mٵ��*
P����Zm���tM@����5Y���g��\�-�>R�6����&��dT �i*7��@���"
.���V_ o���4Y]{FY��������;be�Dbf|==����d�=m�b���U���-�.�
4*׮S\�.�
yM��$?��/�^�{����ϲ�2SGγ����G��d�֯� �H����Ik��#W�BVS������GT7F%yT@g���`̲����R�oA���[r:$�p_��u7����E��� �A��;�'��DA�'�p�\�L�z�cs�p���L���[�k2�lhwhR�Em���d����?Ĭ,�nM�9f�(���-C׺��*f-��5ӑ��xW��(�^����0�S4i�+�N��= ln6|�+�A��*=;؇̊ڥ�\�ڝ>���ɯ�rȉѓ9GQ��ߣ�B�V�O��4<q��Nf��u���sޡ��9S�$��4 %pCA�wE�I@�aB��S?���<��G�e�ךV���~e�H�cD6r�=�y�����%��=0F�n&�f�f��݃a[o�G�懧u�=��p6G�	��ii�CG������w(p~���p�P4�
�����R�~�Go5�gC�#�
	G�Sr�|�	W����l����6mB*�N�N�JbQ���j�y�qv��:�]k���6�3+K�Q��g>,w~\�nb�ZI�
r@���C�5I	�l��S.!�Mzk����U�$f[J'�d����T����n��ە�cT�_3X���v�^�)�M
�6�so[��<|�M�G�S"̕b;P�9`8ף�r�9I�5����+�]������+L����>pU�
��^�m�v w�G5���P��|&8S�bt���s 8�^��U��e:�=�9��(�ۇC��sw?��۴�͖D�������7T�����o�kP��!2���pwy{	8.��ǰ��>y��l��\e~z��}��087r��=r�aK*��)|b\]�1���%��[�j��Cʉ�
	M�'B<I�";�Q��Ҩ9[A��5�mrB/乛y�oQ�g�U�N���K�Y�V/����^$�Nڗ�3D�Y5���S���I��K��^��sc�2���==�o�Y�ak��pL3!jұ|�2�9^�~��݁� :ރ���M�qw?�&��Mh���/�D�{�����&����ܐ����9M⍦���g_���/u��*�?9�hL�h�#�\�?/��5�ZWp���RΣ����ܟc:���q�m���>e��u�3���J5{9��rϑ��ZcBУ-�ۏ7�唄5�o�1����e�Og58�R�'w(G�PP-��0��`է1t��ƭ��@��ħ�*�^_`��`���Z^C��;�È�VN��5�!D ����`�r����4w�`�F�Sp�.��o+6���M���J|*ҟ���YK<j����lr�ަ��C��t�emzȆd8�Op��,`ǌD+�I>{��3�֢"c�p�C����z���F��q���U�K}�7�'��e���EK����ZB#X�^ċ���\m�r�׏�x�o� ��{m��-F��yN��v��ʗ¯����*�l����Z7�9�K�n	��۔1-	z���OgF)�%��j#,��8i�&� =+G]S/36j��^�8���A,�Y�����ZQ��;f�7�Oƈ���;���_zSs�8��o,m��2�9K��I͙�/ND��=��Z^��m��1��.�؆I��8B<����JHQ�����Pո�c-�m|��S��nk�_e�!���do�Jy���"he����JP�r�y 	�&NSf{$��bi
��dx\�*p�0���u8��a�&�籄�m���I�fH��Z�k9�|m_��12��Jl��Z���<�C��)����S"���5t	������WB�[�p����p�}������Z�c�A^i�㓝��z-����Q��(E�y���v�]�x"d�W����<�Ë:����̴������z���В�,����i��;����O��C����wop�! �͘K�67Y-��#Hk����-챙�{��L�Q5Y�U���P��+H*��q>�������U,�(��]�8����$��. ����@��֌�u�^V4��m�54M/��ޑ&og_,d��QI@�^�:���fl����F:�2}/kg�
�-��ط�L�Xp[v��"o�-�
�?V�6^��+��Q-��a�>=�#*Gl���kbT�ԗ���'���/y q��E#��p�x�!1�R��ܬ�*��E�ߘ�H%�,��R]�vVQ`z'ai͵?;#�QM��F]ɚ+�J'r�^��JA�lV	��=r� ��Z��h����b'�S�xH`P��)��i�B�����E��vq�R��+��\�����\�%����	�d����c
 ���09'!(d��B��
�M�,;#�����{%����Jx�u�/K����_<�bC��uuE'��z��S�N�,?!˛Uό����!�V���wã�R�F���cA{��$*������/ssMJW����`Z;��i��``ܔ�4�x��ΐeI"�I,�����;��KԎ���ל9����cä�o�2FMq�+*i��+wKwE$�]��.Q�b�z�;�ۢ?Y�[�gv	����\a�`�*P=� �����i��
c�t|� ��^��"�2����=�f�L����r��!�ch5[̚���jeѼ3�*S�B^{,UMq�]��ʃ�UU�"�u���έ�j�n�i�,|���0NWf�l���pP��fQe[���%V���U�<!b]e�A����G��`����Ћ����?ا^߆u�����V �[Lq�Q�-�\/���]���m�{�������)g�_����>J��e^�7)y�����P�`��v;�4e���I���Q�p�ۏ�7��=���alg��l�+�ہYI�'��7V���w��_�wA�}-�ӭ&#������*�	<��[p\f�렫a�L�?�uC��1B���v���OZ�<j\���QD-��"E�8��^?B�Rۉ�S9��1)�3�9fϩ;J�����"�C�١^~q.	Ι�}k=���tA���ϢN#Xx�bxG��5�x���e�w��u��洊�&]�^EO�����������fI��EI�T9z��N�Dѵ������cg���@Ȯ�b��*��]BQ��}�Z����M���m�H1�.E��Q��ؿ�>.�dޭf�C���	���-s����Z��¾�(`s���M��P|7?����X������=g���`��-x���Kŀ���'�ؕ�/}�+V�fE$.Z����.k��/B(��c�p�!O����x-�E���M���;�B�?���8F��ߑ��� �:�p�8g�mu�����b�j.h�yp���i���\��oN�iaΧp�9�%����.���h4��.CN�y(��f�W���&B�9>ֲ�0�+��S9fwjמ�O^2��w�ϲΜw���r'4�?h+]"��G�$N�Y��Cշ���G������-�������i�雳�A͏��(m�cS�T֟�hi1��ɤH�y�ǃt��s9{�Y�v��C ��k���A�a�֚#Ȭ���Q��%�4A��R9�W���yݍ+�Í�x���gӣ�b�uiq��yA(cx�T�+��@��p��ӯV�I���o�X咵����.�??��_�P��x�Z�k@�O�¥&�Q}�S�}i�� u!h�C?_`#�Y��nQ�ޮ7���Cu<<$����c���R�c�!�F#�j����pBv�����jbZ#KPq{��*���׮I��e�6L�k���,k��
)�*�������ӱ*{rn�+��_�}r;�%�ZK) *��o	M�TE6�`�W�F��Â�!���*�	VͰ<�@EeP���v������?uw�f�Z�B.���\Щ�ߥU}����W2�[�?�r��V�P?����K�L�4u�փ
퓝Rb�J�����$B�<�������ʑa+�7#Q��/h7�t���$X�l-Ծ>�酂�p��>�)��Cn�+ȣ�ZT���Acqy����7���g�L����)��9$��2�ց�KTY[Ocܤ�լ��Z��g��EmP��ws0B@*��Ί�'B�Gu�l	�%k�� ����B���f��k�3�6�nZ���<7��ԕf�W �d\ʄ��,���T�L�F��\&B#���	��T���|.�V���o[�0[@�%=��òv1��}��n����rod��m߮Z�qa�	K�6bg�;���Z��lL�,��^��b�;��*��Y�����w/�u; t��HMGnB��3N�S{�����J��_�bƬ��ج�J��O��!�
c�<l���)�3��J1���Bz�N��/*>Z�,�ǁ6zWm�q��Cd�X��#����B>o=7�nuf���?�Ar"�U�}��_֒�����WzX��o����h"͌p�v��0+X�Ic�wo�{R����Ch[h"Z�a�_�ZM}(YL�k��hn�w�ʻ䒙ũ� &G��+��K*���j+����(��R�x9�;�����.,����j
L�`c~�0/)��c�$��[����i�?���ˎ���X��6��B�Ґ<v��8�w=�p,�)nO-ǩ3$l���-���Ye����]KiNA����8�O��8��"xދ��a��c+OF�#�XO�j\�b��l��:��먜�c0�6.�!��a�y��UͿYEd�&p�3~~����]d�` �, �y/&��#Xl6���K�2�O�#���s�@G�ܗѩ�(���Ȫ�)	�ϯ����q9�:@S�$��1X�֛d�8�+�"7i�G���n��+�咰č��r(e%������9b�d0�,�����۠�*���#l�l�x�'���^pi�(8���Gk����/]?�}6���Us���j~䎑��?3F�z�.�!��;R�z���%
6�nm�N�?6��݉��)r���ǡ��[G�|@���.비 ���T�w�N4�+�L����7U�E��s��h=l� ���7�p��m�������k1/�n�N�Q;�,8����Z*1�u=�a/BMĖ��]}#�
��Y[ �|��K.�����VI�q����	L�%Jm����d�kMXk�B�GD˼Wi�!-��Pʯe0�80�Ļ�S~�&�o���v郐(G驉���Rϝ�V�Gu	TȓBy����/�ҀJ	"WS�dF�TS�.�g_��O�9\Yp9x�y��R2,,7�vF�<a�K���Vo�"M��N��%��_��S�N�2O����ڴ��.����:�0p*�렭�@�b�{� ��%�n���C���y@�A���7T͸ݝ̡�;W-���D4��׋t<�{�,؊�°��]Dq��r>g.���8�G�?��Y�)��1�ˊ9���O21��Ȁ��q+�y�O��p!�L��D���X &��ޚ6���P�%�b�5��gm�p���+0�x0�c�M3m��O�B}E�.�+��>��e���}��` 8�m���V����?���Z��&8-}_B�L4ih��=WSH_�}rR���mI[X�=��ۧ�h�H�\zq�4"����e���oC2ު�m�F��W�}rP51������U������K20���4��fHZ��24���t�Z�# �f�Gj�u�ͅ���:ȯ)M���}��MiS������IR�}09'�q����0�B���Qh�
4��z�~��J�"�j���(/z2J�V��k�lD��9�+%�>���Q?�9�x��Kc�<�� V:2ъ=z���Z㝬��2���To{����jC��!��qkn=rB�AЪ2Ѧ��� Ws"�,_�r�����q�K�s���M���h��%#��3���G�E��c�f�)�<�tR��B��YW����.��C���P��x`���ӷH�]U�MñSW���?��h�+��~=�Ek�W�M<��_
(��V+�A���
��|���L4���g������K�ޫ����%?�<��A�&�{w����?}���E�����A5�ō2�F����KL�}�Q�}���
����a�4�U�%�N>��8��z��w�P�q�R9SX�	�sw�#Rw�o@�����aB�ڗ6�O�˻�Q�i�*���!�-��3G�d��B���'v�ґ�v
Vay����J���hB�hż)?3E]���z��M+wnӳ�c����,hx���F���[�`}���h������%%'w;b����Ͽ����ـ�N��;�5/�`h�h p�$�#T9�yi�����' �[v�Z�v�-�4��ȇ�*Z��_D�|C��-(���;�\��th���q���>o*G��ȶ�C«����\�<���!a_f��y����
��Gz�,�5��8H���
��{�l�!*ƐD0���:Å�Ν�� '�pΤh��VӾ��`���4��[gi9d.�ȓ[�*q��z��Uî@:�iE�B�`@LŴ�8]W �'%}����9�\K(��ko��cù�M͡�����Kzz�趄�[�ŎcT9��Q���Ğҳ=u��8��c��bU��� �W �nCo�C��a���S�[���[%cU�c��fǍ�:���XY&��n�\ �� ��e��b�^'�ke�D�g��4�w�,�n��>��	�_��x�ڳf+�����Ia$�󫣲��ݺ#h�:�C�%zA�|�Z�6kC�)��T�̀�N��W���>���sX�[ �����8�<6�K�^��/��3���mفf|�SY��N��fi�2z	�ǝI"�G�Z"l�	%�;��%�]�$��Y��$k�OKJ~D�B�Z�r���Z���`2�5Ԑ���\	���@�<�1;P3&�AITVPw��44߷���Xg�e[��z�X;�}��
��=k+�͊�yς�����p���΋{���y�hu���Q�D1��C6N�D�u��12�!Ҋ��A�M�;�������~��Ќ�\�eLh���'��?/9
u3#�e8���#+�H��"�':i�~�U��mdg�P���3��@7�7ރ��a�H}��A֕T�@A@��U�i�P���=ה��J̻a���0r>�SL9���F�r�g�
`\�GA|�o��H�g]� ����\��NG�k��а4B&\�ٯPa�w�1}��<�*���%�s>�0 �!�L�1m������a�U��X�$����bDeʆYV��!n�����e��O�+�����]K�B�d��c��q�]�����<����r���Kk� c��\�RD�D���`7X���p)6��n�9�	�V�e���Y=�y��?x~��u%���J�ǈ�l�5�+|��6�`'���ޑ�Ns�����I�G"�@��&����3k�up�{��6�J8�Ș���;p���Jΰ�:v3n�F��ee�� WCR�K��̺��Sro��MU�Qt8��@¿;mE?��P�3��-�`Mq"�r�1����"��)@���	�.4�)��t �S����,�{�>�y���ճ(�3k��5��� ����A��x��F�(O�\B�c�}�B�>4/y��3�y�;�%FUjJ���T����f"�>����W��n�\���XnJ�W�+V�&�],D{��ڥ3j�	��	`�Y���w'3/KQ=L$Q;�g@k��J.�uEx��@�*�FZo$�EA�O@O����������$��w�{�$�K�P��]��5��i�l�Ľ�� y�&�!���O&D�S�.�QTȶ&uȯ~��{�f�S��[���X���TIOϨ 9�j޾J�]�z�V'���b�:l�H�v��;	�DT��u��~�Q?���0���c54�0��i�u~�'�P��x
1?���5���w�T�6�j�86�(��-��X���l�RE�l��	��/�	�N�+I��˭Y+Ϻ/���g���Ř��D�$Q�?�\%c���of#�nW�A���j���W�dS��#��V���`��_PK�2r؆�X�c}�GYG�3�:��~rGy񈿐�k�86������b7C�jy�	��X�ϝ�p�w�:�9�ܺ>���ElG-��-��`v {�tL'�C#��^&T�1���5�H��Uܗ8E��w7sW��C1\����C� �lP;���?$'��	����^����NP�,\��St�ES鼂z�"��ӇՈ��Nϙ4�~�Ӑl�@(���bPl��AE�b�Ha ��) D���p��EiE�5���&A�Qo��*�O���ߍ�.R���z��G"��U1�)�����y}X_�U-Y;�P��X��I�R��Ѷ|b�����ķf������UsxU�L.�XlW�e"Qd�s
^d��ݥ�޳���f�����]��Xs=��(t�S�+�'��hPoú,?�}����}�C�iV�ۍ����1��o�{�f��ɸ������(~T�WpziD�y2�!a����t�c3��'��Y�'�ԳM5$��R�iR?;=C��]�w*LS��K�]� �j��}�ô�v��sq��.�䋋Jh��(��n�/Fq�z����zw��25ӗh�U�Z���u���<uj���&H�T�0m��������g�]_�Q�����3{t-�������X�p�Yc��}7� �(�l�
cTCȼ��.�I�lu��̸�����kz��_�_��Ump(J�`�S�?�<0X��O+����e/N#򨨿V4'��O�2O�� ���d���l�M P������_D�������3��\�@Z�|�1�ed����l�'ƊEd�]2����ZV��8���nS�t�t6t�/��N.�֟�X#��_�i*+��VJ�"�n)�j%�)s�d�$$0�<���x�@r�Vԕ٭�U���D��;�4��(�y��덠����:v�x 8m��W��0!~�q�:{��lJ�E�����g���;9׋�����.OX;�8}H�_3�Xm���˻n�^D�0�s�N�x�S3�$�X��O�C�hrL��~d�m��T�֡xfo�;�E�`�����2>�Vm��X���"�]�+X�W�nA�HC�>�P���b�3~T��9�Y�uC�9�,�8l��x�w\&���[��|+ߔ������&�e1&(���VuH��\�1��̲�M��
u7�6�'�$��`����ѐw�+x�YoY�)�x�Z�{��ܷN؍<E���F�l����|n��0q/R6t���mu�(���z�A)�]
��Hӝz��E1]J����N�X]� �����a�	�$�i��L�ޕ	�_��3Ǭ�ҪX�?Dfv�d{FU�!�(�� ve�EP��@�O����*[��Ic^���|������&%�G���|���U6���`Φ��p2L����X�n~��^�m����i=�P��+�ُlyp��K��BL���PA�vN� ����v����:~�F���fD?�RP�$��}�zgx��t�	� ��P�҆�T]�߇����"F2�o�Ш�$e�Օ�X�`*9���v��Ȗt��w���P���SA��[=���f[dNTiK3rE��/���I"�I�� ]�M��mDJ�+UGT�n�9�;Q[�C���▦�-�m0���O���m�S�ݷƞʋ��ї�bD~�g_��%��c�s��T.C�-E���B���+�n�e����A�gN��f������r�ۤ�Z�����Ax���S�_�.B�Vѧ�:�G2���y�(�x��tY�/A|��Z���ȳ�d]c�V�]b��L�Z�uM�@SlP�z�Vf�c�b��:�d})�{ ���@H�6i���8�q�D�1;�>9�#�ۊbc�i4t��J�c0�k:���;{#!��m���]��_��
��+����\��f^����J��nsme�`^����a��1.U��H��\���eK�8g���Eĉc�uI`a�lS�( ����(���w\Hէ���&�gL
<3Ɏeg�Y��K�Cn�A�����i�pc���x`1@W�ʇ�
�lY�9��mgZ����j�I� 5��)����0�g�W���ܸ�JA�v�}��?^RҠ��e��=Ez����_���;� �����`�m=�~i8��DzX����{�b�S�ٷN��p�_���������v���ثaQ�Պ!햹��Ò�.�.�?X�h��j|���d���Ls��Ѽ01���1&����yCWj��n�������2��L�,��q[e��\�? l����`��8���.yZ��#�|�g.����	�r؜�g�)Jz=���C3�?}{�5Vܶå�2H�!a��p�����sM�O��hZ��b��'\�����/���
���ԧ�X�x���Z���2���K�B���]�"��
�5�n=5����:���';�+>�w�3���V�llP[r��FW6��(N��1;W����v��<K�HiDQR<E�v�s���5��퀩[^A�ȴ����-�i�x�d݊�� 4�6�y��:ُ��>�RK8���~�b���}�,t���+�����u6Y¸�
'_��ծʊ�Z'.�C"[֛���dҬg饈Mn����ڟH�!�5~�Q�]ۭLl�Y;��-i&˫�������zb��Cقe?>{|%P-��_=���R�\�:a��$����J��l&k�݀�l�f�ډƗn6����-� n��v��=�3\w/d��a�v
l/|uh�4�('`t��%�0{�o���Ru@e�;|�ߞ��L�\��-�v���B�X�]*�"m����j��[; ���0�cw�q�a��3�c��*f���'�V5�,U�O��j� ��k�U�iC�)�a�Uz��=i��ݷ��Xs=�,-z7 �}�v���?��3��7��2�*~X�"�n��A�<%�+����FF�$0-�}��E�c{�%�qo΋JD�x�C�~�)�	}h5�$T��ձ)��3Kv��(���f�P����$Q}/q
~�ľ�pYW�rt�S$�9?t�-�� 9*�y�U�����g���
(��|��=zg��"g>j��;<��2�_Eř��܋�U�e�5t���u�R	��=n�% �F=6�d��Ϙ?�`%Z��ix�3���]5P��<f�.Ĝ�u�I+1Zx[�1��r�0P�#�V�ܝ�ҩ$(�+ɭ����̶���'R�SHj�[:�@�*9�w��a�wm.ݎzD�#?�o�Ua�k�J9O��z�i?�M)����zY��+�����?y��-���1-�>�6.6��-��S�#"EN L5�
�U,�H�ڽ������&�'���!o6�]:Σ������B���]�D_kgI�m�z ����U�c��V}H~'�K�H�VyL�l)�i���P�4w�3�y+t�1Pp#fޕ�j��/��-`E:�YϟyO[~2|��;�x|+�1�(�GjHG��QQ~r�w;j�}�b���y��0�T��5��R06X9ٳy�]O�"����o9u��=����wW7Xɧdtlx��gm:���n�iio�'�?�q���N:k�¢�x^8�@C+,<���b����$�4[[�%|�+��xeQC�ݨH��`�Փ��vI΁�����[��ްډ��u�C�9~Z�
��'���} KP#�B��3�il��g�7�y#�τ\���7��n@m�(�~��
 3����n���ݰ�/V�pQ�w��/p���ӕ`�t�fK�"� ��2��+��j>C'��n�.�c�I�[T�=6U�� ��� x�Q��'�&�ֹ����9(��I"~����$Q�sʭM�R;jOpI��M\8W���/�y*CE<�h��X/E�o�oT���F�W�4�q��;l�o�i����=��36�0.��h��Rȷ=k�:I/��X<{� c�.l��~K�EΌ>��F��U��^һr/�Z�ߡ�#�EA�O!����k���N��-c�-�x,�Y�B��z�]n�{a��ߩGӢ�2\�8�y#O��������m�J�%ܚZ�5��$���-�ؑ��4##��1��Rn�ʒ��k{	�P�!MC���!ɢ������4:|`X0Eh�b|�o���x_4]�!�1ݔ$/�/%�95H��oy���4`=\w:'X�/@ڳ���U�T[Y�!.����B���;�Gю�� �I��&o���w>m���W�$�7�1��jP���!�+�؜w	�������L���:'mB\ Y��M�PMEiĐ�ț��-���W`��7JQ�>���ވt%3�"PUk�$B����]�@ϩ��W\�y��z�G[����1�壕GAr�=�w��*��~�lu�T-��M/�|YAɻ�.X9҂&�|�4p��ӣF�����6��� �a�"��<ݑ�UD䲖�2.���1�gͨ7A�ON��*+�K,���-ƈ�RQ(�;�<������Z�.�Xq�ѿ��Y�37���8�8)��� +][/<Jc?���).S��m��N��4�[���5�ͭ���Z1$���Eh|^6��
����l�sR��.����R����z7F�D�����k���,�u�����%�	�ƍl�Y}nW(�tZ��X��tI����s��C[�$�fp�#?�E%Ŧux>r��f ')b�\��[�s����9�L8E'�WԢ�!C�aէ�+x���VV%����b����H	��Pj���3��Xl�"u*X���'��J�<�kAAz���V�a�ԃw��i���f��ajQ��tj3��X�ƹi�a!ep�_�L���*���B�k8܈+m^"��W��6����&!�[�HL�p�5K�X/u/��Ο� ͣѰ���ޛ[V|�Q����\|x�s�-O��+�����	\'���\��	T{�ױ�j'��wm:��[�~�9�O������w����}&���{�Fl��J�y竖����U��*-m0`�$f}�1U���>���^��A�MϤ5���]4�Y��,��x,@�d���)���r�=��$�F�`��#�W��Sg��f��������H��`�4H��H*�3��C��)�x,��30ɉ�.b��vś�xl��cbm	�2�����e���L��v"ڌ�9���V���\7h�t?9Sv�k��Y�ҥq^��ڮ"+�+٢�XCa�6��q���� �e��W�����HH�B��j� O���li+��J��)�i�������I��1��W.0#Uq��r�Y-�)D>ZP���y"ڙ��ɸ&���C���B�l��X�͵�A�������;h�����\�p��)�[�z�mn�NN��z�ؙ:l�?j{�c���xV��c7�滂̩�w�� ���I�_�@�=1)yWLv�>D�w�(�P%����]�3#�e`Fw+[�"�i�ד�c�^lb�2�~> �,T����R'�P����~��A�����Eʗ�{�^����K��8uo]p1���YA����Q
��%#�0��'�ʑs����ӯA{b��Ǜ����%Ǘ;H��r:wL�2am��9��y�PgkStqSp#$ls���ٖ�H�՟h�v��Q�b�_��ۍS��@QO=�����М+D�P�r��:�~�X|:�br�	����c��&`����fգ�,b���c����"Cu�P1��)�ʝ��9<�V���]�:1����j��5)lv��W0
�pM�W�G�&�[�T�Ħ�B�1���S��ﬠ����Z\ЌP���'Sd�E%*�b�|����/NJ�g&}.n������������M��g:���C���ϝT%�c���5w\�*Ӳ1�ˁ�Hkx�;³ј�!c=��K�J
c�Z�Tc�͗k8�`� �w�`��_g�x�+�6ܿ�����l�08�Z��?��S��%+�Ǖz���o�G,�i�Xd{P!��p��U�"�4H��e�'��I��5p��x`���3�X���R�KT�����!R/K�V'F<�"3,��/���=r��n��:u�m�����[�� 4��]���!�ܴ�N?��0��iV1/k��;\�`���qV����B���J'��_;�-d��jDk'`�@ڗn_!l�U���
����{���g����mu8ӛ�&��F�����Ϧ��騉�����*O�gf�l
� _�t��_�Μ��H�5&��-N�����o�5�k�$�4�Gͱ=i��t�,���YAK�O�TB��E���a�n��4����&���"4�*��,w]�>���fh�KӀ��q�~X�x�`|;Vw,��_�T��VߕЮ8���+�-ĭ�g����>۾��j��������\�T!(j�: �%�s*�YX���u��?�;>l���4R`V��7���[�um�Q )9�]�;�^�-��s_k��z�p��겜.���Ĳu�n��D��)�ܼGs�cJ��an_Alήh��QR�g:�L��Ģ[6��d��h?y3�����i��X���?z��g]C��=�bWkj�V8Iq/�.������*r�ndܑ�6��:�T�k�x��������cT��s�*K����9+�\O�o@l�0�R<�m�g'$v��ʆάzP�<�K�|M�$�+o��^�H�i��h)���s�}4�c���oPD���������P/E����H���#��=�r���0(�ܙz�F�&���B;iw�/ .y�Qa8��iH�(��,5Uh������̡4�N�*c�*�'YʽrA��U��ۚ����ŏ(��7ָ�c�ݾOY��#���eUT�c��	�坋z���ɋ�B�wU�1cm���J�@/�2oo2����6{�;��/�E�7���m�)�	V�\X>���
{8���.���� �O�����[[ŗ��� ��?����t;��A���(����k�����=2�Ncߩb��NIo'%!?SF��w��g��.%y
M�u!}�l�Tj�
��,�qhl��M�l�ѨN�*��d�c`��,�g��8_�
P�:���:_4k���B� k�Ђ�I�Ĕ��i�oD}��&:�p�qj5,�c�&�SN9՛����^�2�_�+��㍷?�O/�]����	�Y�K0v��� fnB�e�`�Ĝ���Nf{|��2#5�d;���ѻ������/L�n]z��k�=�J�Ͱ��o�{�W�jk{ N����7�_t� ���e�$SƸ��^t\J�~�@Z6���M���]�FU)o
A���M�H��׊�bLU�������&l��m�n�kև��H�i��<�6n��W��?g�B�ZΈ�s�^l+��Y363��5��C���W�Xݍz��j�O�������+x���O����˦+�g��p��u��y�΄�"Zf��Oĭ�p�}�C6�n���Ӎ���_������(2��w�B�^�+�B��ݑ�T�<�ˆ����^���qL��[�:*�m��?,s����n>�ڽő�1?������J�8ݙ�(؋���\ۯg�D�oxJp�I4���gx)`Ψ��7CD��;�X �ɋ�@9�Х'����(Ϣ�7�/-�� ֩;� M��K��}��u��I�����}�t<u"L������=���^g���㘾��a�,��̽�T�\y����}Pm�S�����Z�[�"��W��,?�>���+"mc*V�8!���MZg����K�G���H�>�*_����c�҆c��(���&B���<K$��K�ڔ��������H 
�/�D�����?hJ��� D&"�*C�C\������V���}��T����ݫ�}�@0;�!��ѱ�W�3Ƃ7'���Q�4�Pxs���o�r��IT��ft��!��`� Jr����x�
jYET����C�SV��AzPFɣ��Gi�
�� BIw�k˜�/y�9PO�yGs�ݱs���:�"�nX38G͋�h��u�tn��OL���3��ӄ��1�CO�����+��Z�O��ME���(5�0G�"�Y�~*�#�*ʮƀ���[��wg-�
ۍ��L��沕��n�1>�1M[�	��s�����T+���M�?�)��@���!Vk,m�v���U���j����ҫX$�V��s$������.�'aq2���o8Л����Bqi�w%���~gNi�/͗O��>D+�e�O�ؿ.��/�	�iĪ^�������C�j܂K��J	t��;�Ne�So�E	�C1�r�s�:��
�I�5"/�S)�@��"3����#
����G�H���}����<X�X�UL��p���j��g2I�O*!�\�!��ޟ�{��[=�MH�� ���z���u�MX'��0j���A��:W4J.�&�ð���,�+��4��Q��������g�Z������q���ML�i���K{,F��E'�`BGݕ<~
����@Usb7wYkhr0��u� !�/�E�g�9����Ɗb[��7�BR��d��-s<���/L	K�;W��??��:�t��pjY)�.v�\�:�[C���,��J.oͣ�*�BY�Ғ�/�mˠk��B��%v ��և��u��@����c�M�b^�C)�����q(�,����%�t E�z끞��ٷ�u�U'K�S�L5 ��@y�e]'�c�t��S6��aD�M�l}ͥ�5:�����=��Kn��{�<�{4L0o�礟QFq�����b��z�J�h��#���c��������x�
�������x[���N,k�x.�y��c�G ʎ�z�L �� �S���`����Ν	e)emRp&��'� �7NhځP�*n�bvC�4�<M^�;�
����K���`U5�����I.Y��Π�����`H.W,��;�|65��Ly?�O��8&At�Qף9�N���H�z����͒d�U��� ����C���M���)����
fTYv����� %Kh���>�:���o���I ֕۰�rK��@z(h�?*�������H��"��<w���� ���VV��wb�Ȋ����s׹�t:�K�������]�\V�>���?v�kT�j�?R�${�@�
��%�2Np���}.3H�=���eA�H����}I��J�n8�쥣F��I��(��w 6[�:��S��R�Ec����lUl��f�8���U!���!�IUㄢ�
����o�|�43�n+��i4&Bf��n'�V8�N]Q�MY�FÛ6w\�JxtZ����LnnZ���֘�f�u�V���}�(�| �ZQ5_�P�@��K��U�)[K{��N���,��
d��*���%�"G�!1��+4�11�2�������q��G�P�"���*\�����Me������w�D��[H�1.>��Ⱥ�ʙO�m]�������9���OmD���٧�PX�U����9a���7mzGG;�d꘭��W�b�
GL��R�{��
�����*�W��J�����{4� {������a��d�e@�xt���e��ivUW���ھ��s��.fV�g%���%j������хBm��p��- wR,�{i*ʔ��?!����gz�g Պ;_�m� ��L ��1��-�W��X��֬ƒ�z���(^��ib���co��Iܣ����y�P47� ����s���SMk�=��J���c{I���ݫ��rd<�	�����p^����y(�?���m4q��0�E>D1��c4�| �`������Z��Y��� K�A�$��0L���jW*�Vϸ��ϸ�,�Pv���B��*�d}��I��\�P�>�b��l!�� �����N*c������SZR��s�W����m���K�D�o���}a��o�j�T���ш��4�7��q$}���R㋨��7��
Gl�`k�$w˨�ӖJ��yg
�oN�۞u�ֈ%K�N�(~�V� b��&o��Fϐ�k�Q��T+7�Ѫ�,ƺ(�븶�v�	�������Z�ST�O��_=��`. @��4rt�-s�=p֨URr�t	�Ӆi�A�v��a�r����qjͅ�S�\)#�@6Hu#�77P�w��_���m�I��g��u���p�%�q���,D(�]��O����Ip�ݝ.�<�}*�-��9bS5�zD�CZ�>|힛��G������k�m��a8>��0�S�fO�i�e|q��)�.�Ob�Ge�\�
"zwʲ4�H����x�H����r��v��c�@�%����Ph>��}<��xnT;��_���7��N\"9
Q>c�l�b��4Os�x,r�_��(f� ��(?��jl���q���r�R-CIM �c��eu�v�Z�u�)]����&�&w��n��q���HGD��H�$����b.i~����N�ȇ��FNȇ�&B���i���Z��Lkh���Ց������G���>��yY������CJ*(�L=)T;���՞���d(m+ñsQ{H�J
�q����'@��>U2��-ƵA�T�kKfoE%d���y,?MP8I�r���YW���<�*I�䁧�dc�9��٤����\��$���wR���Ե�'�ND`	�pTM)���ٖ�GF��J�LL��̜� T�GA���⫃�!՛��u&��3L����Pa�Pʡv/V���fN	�G:����q�K|pO׋�uƓ�w�y4�	D5��<���Gr1>�D��ߣpwd�k����Z]����|DC/�9�����~�ܦ������~-|��Fe���1���螇ӫ,�g�1�.�cqOf1_AG������/%�j��*b��N�D��} �ܓ+��y�xG���ߔ:�:��Zw�R������X��G�����Z�wW}_�+��+W�GOލ"٢��+�f;W�$My��	��{���������f���s38��'�&8�?EQ@�BH���CmIn��+��eKA`p' � 
�d����x$������б�"����C��D��x՜UV��1�c��GqJm����<���zz����������:�'�0QNCxnp-����w�@���g���ہ+���Z������5����>e�@}w�{#a3������S,?wU���[�S����i��� �	�n����Xe�(i�{U�E�wd�/�S�|�1�j&��b�-�� �0翻(@5z+sse�(#�
D#/�!��E�����?
"�y�F��8YP���S��p�����%�_Rm��,��ʃ�v��Ԓ-��X��%L�B��U�ǖX�8-�K���jK-���*O�v���VR
���.�Z&gi�R��d��H�z����R��.��do�&���è�s�.���n�I�.��m�5C��yM��=���	"�Y�x��A�&�hx��Z����b�fG2 �p��]�2�>8�1F��,���~ �8�*I1?�<��-�K�V}�5����)���I�㔹�g�@ewfV`���B{p96�ݰꮑ�4Tfj�-ꇍTY���P!zXji[�a`?0��������WS��K�J'�K�
��[{�O&m}�n�RU�x�t�AI,�1��~�U.����i��������V%���]8eP�i�lH�K���Dÿ��i��]��c8�~�L�+�i��D�-�JR:��m\����� nv��x��-�>�)2\~���x�������T�avw6�\�ٺ�G�v�()�y�������I�o! �.�����zl����Mԍ��P#WͅCT<P���H95.0�`Ƞs;Tk�̂�=�1'lyz�R�aV�!z�!���\���C�mGPU-j;E�
��P�`��dq��؀�TA���ڀ��@>g�)�X&�z����}��/C:���t�A�u&���2�c����L�?+-���oT�����IK%�e��T�FO�����Ǟl�a�*lj�2��7��0�sb/�}v p[��.&X"��HSl3��4�5Q�Cui�j� �tyPV�1qڼQ���!q�
&���M�<��}�Mpn]:�/I��O$�i��j�ɡ$�mT "]/�]!�a�dQ�*K���V�m �!���}:�V�Kq�8x�q�qnHk`�E�Y�y\.N�ȹ���ݗ	[�|J����޴	��w�#%h�c�o3�MG��Al��JW�/4v�����n>���E%��%^ڗOpd����4��U��i.��C8?64��o8F"{y�L���i����݂=��o�$?�3��6�vLC�A�5Y�HA���&�P �	�BQT�&��Q[AH�y%zX��8@U�dM���p��k�n_{rS0�����D���\QM�p����Sq��"������\�0�+��J#����wԞЅ���L�l�]����������&�V��v���
ix�ΰ����8@#����3��b�����1��j!����r[j�u�����:h2r��a������
yS�+�\0� b�н0�Ѹ����o����O���?K#��<�?�?B�"�?�?��ǒNnr���-�e_ ��^b�H����Ӱַs�S&������O��%�M
�����t��:��u�L����@�n=O����s<����_/Y�]4p�F�������0t�1T��рR�P�I��`9�$\(n�/���	v���x~��%�L�	�g1e��OEm��ytΒ�z���2�t�ؐnRi��_�_�H|��o[L̊�3�!�x��l>X$w�0m��t�\xj�>n=�����T��͈@��;y4����B��@�kt;�c�������*�v��0,m�Mu�֍w�8��b�(Wڿ �޼s���m����k֍X��v�Е+%��m�%�'��.�QC�����9Ыq_@_���=gCO' y�B܊��iy�����}K=U!ӱ�
��z/?G�p�!�W�Q^���2R��KR(��G�#3$יx�u� ,��u�\�����ޖ=�d��
�o��m�W��X܀oge"a�K�w�@�E2�S)*l��ɺ��53�Q��?TP�ܯ�y�OУ�(.+q��Ad[�J��@V$~�)�OXj.��1-���$R۷��k����ݤ1�I�W��6������=�Ҏ�9�-����3��R���|/�Dq���k�
���_{w�dSX��]�&����P�Vcoď���G���+h_���7�C�}�8wd<�:�n2w���Ԑ:��bu���Z8�B����v��Iؚ+-��P�����,��_r�ԟ�g��tv��S��G�<��1�8�#ZJJA�y*�������'7U�E���=�"�f�Ij\�&�� !��+��ҜD�(���vB*���<���d�����l��U���g����
����:����K�%���ܜi��@��X�RMT&��%�Z`�S�_M�-�w�
�h�W�mgc�D��d�����O��rP�x�I��o?��pH�[��J��F�%��#�,��-�|�w��*��3ܬq�h"�!'{/Eh��-YZ�G�+Nt�������E`������f7v̖�o/���;�@~f���5ڭ��M@]N�<\-�N��[%z ��N�m|)ԚQ\��=����^t�8 ���������:v��е_�b,�;�����.�N�:=�&�b��lc%��b _I���(o��F�����H��D{k��Ns4�2�a��,s
<}�iw��52p��FMM)�T�E�QB�%�DK�(�����Q�Yh&s�G���]_���f��"��`��ր��q��է��}��E�n��Kv��o�r�rDt͹��+�~��C�C4ٯ�k%�B��8��%�׫��;�K�5�#p��%2�v�8��W�aj�2�(�hわ�<�q���y���V� ��qt)�����yd�����%��
�����w��0�З�|bu�F囙�����ǃ��PJ����K���@�%��'2L�(I�5���4}��s�&I����6Vh!�p��:}�o�>��iem�xmq���V��j��D��!�H?��앭�l\���p�ǗCWQ)�.�\Qth5�zps��R=T�+&��%nF�_��?iqف?������I�}�-�9��eC�Bf�J�
yt&�!�⦛AL�R��⌉���.��1:�+�A�<X"7��=c@f^Nc�.i�c���d�ްTGR̵�Д!|���4���3�B݁����n�9�g�ܩ��4�����L�i��FC��;�qr`I!o�ѽ9���.�"zP�g2�����=�b	2�4��e�Ȼ,e=��{�n���ѣ`t��m�|��?ڎ�~�����X���!o��0H��Rd�<!����P��[�*���Q5�#+a���`��kAޑ���W��7��7�� �׻��K�Fo�o��СB02�3��p�ﯥ��4���s�"\l�!���У��
�PT��B�"",{$n���_˿c\x�oELr`O��;N`��̥Cy��_^�:G���g�3�k�ֶ���l�y�c�P��`vo�)���7�]󃥘��h���_�-���k��`��S�\�W��-�W��.k�@>໳����:����i�V�٦'yF�ÿ�r�����Tk��!8��z�9g'�-<�G��R���.�yrؒ%NH���������l�5���=/�/�~�����G�
�-c+���7��R�%[T'υ�E=��y��_/b��O,�}�D�UҁwKj�⤇<ؕ	��[B�o��\�N�/vy�����P�Q-[�j~��,|hJ�K6�1��yfC	%�`�,��M��L��4]d�V�<[h��]_s���n��?������ܬ��� ܲL�6r���_q��9�9����Al�&�Қ�+���b�#S
��u���(�sn\�'/���� Vsc`��жm�>�p󌰠�?�"���R��Y���]P�R���C�Gf!e#�*�=񖶃�J/B) 3]�Y�t��������xC�� �����{���m/�[^m�M��;R�T0>~���4���ht�s1X�G�E���-9S��wW���	��6�֜�)��ݾ�M�{�i�}ufkW�0�8Pdv%�3>�
>�J<���V�>iH�c8�ϳɤ��� ���	����������o~׿�$�z��yA��m���G4��`?`<�P鼧+�ۗ��͘����{w,X����(�@�6a�a���I8�?����2j�^�.�o.
i�
�d4h{���ꫝ���E�K����هs�+�8geH��~YC��$����滅`�ت�`�DBʉ�#���mb_MJR����#��bX�Ξ�9�����q$�d
�O��'��_�ߐ7�A�σr^k7\��1Ton�L;;�ؼ<}�1�\�ɘ���|�0z�'�F`�4..7c�s"�v�'s�b�^)��D�*���Q��<h�C�I����x����E{	�r|�']���*t� ��G���2�N�]��w0F���!�wV
xf�_����.����uqx'�0�ǥ��@�|��3ż�����AEhw��*��DI��s��"�uI�,�\J��%�?�LZ�B����X�1U�u�?0���,t~3�0K��A�Y�I�a$�_Ht�41���i���N����,��Ůe3�Z�^2l��s��P�ܱ�~g��|0��Y��:ݫ�b�}�Zy.y)�d
?ܹ�[���;��q��vO�%�2����Q��0�ܽ�/s�V"r�ya���`T��b�X��+��B����yt�9ﾶ��R1�JD�&��P�]�Vc!���bӊ�l�_�i��S����ĳ	i���C6�q甫o�u����7�,C�kLYOxPל�d��J�w7�� �Gm��cqI^O�ܢ�@x�W���T/���M��U�wg���	74���S��C6����ݶlDm�9�y͡ID��?Eǎ8�;�G�4��+k!$���<�T<�SL�4Sq����>���| ����	/~�<8o<�d@�.A�>k�s��}�FY*��:tnop�B!tzSV��l��D�ɮ��v�β,R_-�b�d[^�����R�8�I9ī�\uYS��k��jxjA�R/�H+ �T=j+��4�!�I���H�6�)1�����U?�ђݙ���	���7��t9�����r�>��'�Ԙ��c��T0l��ׁȷ��z�VN�1j�X�t�ހE0~����'�u~ˣ��N>Ħ"0E����ty����V��p]��7��g��K/5�f����~��E��l��%`.���������)��(F�?��t�9�`�c>�������p푹����?�����y���dAwR$)�o*'|�5,d$�DZE��{�Q��t�a�мB@�i��3��r�Q},��Sf�,�{��mq��t,�n����KSJH�O�VJ�Q;��$GK*@�<��VL�_M[���L�g9�ubVo�pHx`��:�����-�bN����e06��^0��L�@��]�h��vZ4�+&׹��1t=O� ���k���k�w�jE!���_I�.)�g�ê�Ŋ�j�a��z�s�p��D�S�l,/���,�G���)4�(�L�-��;s���9+ZN�a�e�փ���g��"_>�&7�v�~�kHt����t���[3[uKH�MT�L(`���:��}�{�v�b�,�#��ۮ��g��4��E}�P�XY�
����/42�ko�=���K���/b#���J��L|�d���D���p�����������x�-�g����YvFu�
�~��i�Zh�E`|'�!� ��Lg�G������3�O�鲢�Ts���s�c��t!ٿ�/f����y�����{��c����`��s°�Y($��$񋅨:TM9�n	��J��$�.�"���!Ǵ��7����ss��n��'�N)�k�	�1�b\j�4�8�~���B��Bz��a�������D������!Z���� �?I��+�>4r�=84x9L��]��ݓ�	������!�����OM�����;�*�S�C4�:#��-:cQ��)q�@E��ϸ53ބ��D�V	��A��a�"�=�㛕
���c�9yR��F��+_Ct�U��zd�^�e�Է<�%�AW<���L�����t��K`�=����iJ ��g���'�R΄7�q�֑���(�_�g��s�	6��F���z������j̤��>U�!���[���D)%��P��v�JIt�����/�����;�����Cl�
������2��f�f��ғ/�bi��y�J9`�>l֥D���^�`'�?�����й���ɥх7ɷ��:���Ǿa��n���}8��+g�f)O��>y�,>��[��!1B�l��Q��k�yJT^YfG]���Y32���&Pa3��R�g���lց>��Is �����-�es��tAB+vƟ�}楑`wܘ�.�p�֓�7,A�w��J��d�������s�%H̟��hZ��� ���8��KQ�	z�H��[��G�$znҲ�����)\̈́��rۘ:���&����I�?v؈^�;;��p��?D��&C�		
�8|$��:^ ��ŗk語qT�����$Sp5��l�ܾʙ�ӜO��P-��k^�������,|��PL`ʁ}JV�A=���`�%!�OwWY*��i�&)��v]bS%���kFB�S(]��~.�Ά�3�;�4��+�W�}�Zb�7qiA��5��J��?.Sk��7�@�@�#�WN�b�~4����2t���J��0���O1��R�>��Pƈ`߂�ւ��v=��-W�+�q3��g{.�����Ba3 ������:K�[OJ��C��,`����M	d��V>�-�X���9
��0��6���m�s����fq԰e�����R�=�Peڼ�V��X\�#��5ų���T���?V�!��xkO��3i�$d��=����E�/B��]T'F���]��S���|��m�S�7B�j�u��H+�7y#�:�L�T���S��s��J�3���d~W��'c������p�,VF����=�h_܄�G���MV�~�Pq~��Ɩ7coI[�ה{��}v�j��r[t	��������&}"��O��3����}p�p�C�dp�x&���evI�)k�]�,ֳ���_�ስ�M�����p��$�B�j�����ϖ�-%��tD�����,���� 0 �d(�\���� �f�E�d��	!s�:���+�dާʇ�.�)��ƊC�XW���#�o"xa��c!�g���i4��ѡF�u�6�L�꩘x&��)Q�t�a�󜡾��IwE[@�3`)���Vh�N�҂��l���	�]駏�F����s���h�9wUՎ4�	��tys�{�Z�W:V|B�A�a«���:��B},��Ԙ^� <���}|��շ�=,�9��~]��|(�~�/�oIL���������+J&yo^=Ro�u�t}e�,/�d����/3�Ο@A���$;hS8����9:�` 7�ã�0l'âО�o,�Ȓ��	V���4�f���0�9��|��*3�#U�3�`&�//�
�!Oh;!P��)�/k�{�����G��\�}�-�P�dJ�7�<�q���6�6����J���#
da;��\�[-Y1���ct���9���
�a���1�:	\m�@��~���T2�A��6l�Ju���	j�T����*� �Z_�N~�eTP>�9�n�F�9!t��x)I� |y�i��(}��M��/��LF��E��{�M�_��͐Z[Drr���)��u�h�QE�S(;�v188*�eP�=&�m�
�.�(}���?8��i��\X�����?�d�d�VTW�������DY�@�ܺ$��1�\������,_�̟�r����s4vK���U&����& ػ\�Af�����x1"����j�W�hW��	 �\������X{^�>�7E<�7�2��e#����
(]Ǡ�ƀ{c<�F�n.�v2�1/|�/�Ӆ�����u�3�Yag��[�w�[ޚ.�P�J�=��|�螇�3�� �8����|ʞ"���"�1��d����V��J�?��-���"�{3~�Q��dA8�~�M������E<�\߬�ٍ�����5�XK7�@�H���G{�T����	h;H�{��`��e+<����!���u�����4I�����Sw���������کi��X�9�l|M��ۛ݋��I1�0r�JY�� O�H��J}�UmvR�Il�;`*A�3�~}���M��KE� CM5e-ý?�J�� ��W�z4�h1�x
�'�§�L��=�#�w-~�����Xn&.)@lf,N�O>�;%���/�K�aT�ĉ����mz�;܃*Ezp˞�$�'��� �Ш支��g7�D��E,R�.#��V�;k7�fP����m���U�D+ʇ��d��P�GkCw�/�h�y
K�*Yt��-���QV��?~�T����dKa9��XCaR�O0�Y���|�p�/|.�B[��]��N[ ��Ŷ�܈u��}�,�К}�1-�i��&$���%-s�����++wy+R�.�i��g��䯮��ã������	zݓ�Z?+(��a��;nw4�D�;5C���2�>5B&�=��\�L��s�7>�wB�����;"e�..�����6[l7ͽhqo�9.@�X��Q��5T幮Ht�b���.��뗸���Η��{Dg�	�_��e� �����$�[���h_�j�xjp^���G��Uv#Q]�dw���V�17���t�hGQ'������|���L�T�PB��������U҅�J�!�M����)�r�U_�:W����\IV�ꑚ,)뒬�֜�K��rQ��{FF�����
���s���)X�mL�0�Bi�94�u��~��LM #����#*
�Y�����L�"�`�G��;Ġ�������lJ���~kF����ܢ���_��<�����N�ϙ��1P{����d��èA٢�b�����X'V_�9F���y�";��a>�R�b?���'h���\�-Wz
�YZ���l�����F��*��k�;C?y/�s��I��o��_D��2������T����R�4z�=S�ɚj��+P��K��N[��%4eC��1�H��=�3�m&��+������a����u,Tb�p�ێ;��> ׼I�P}��K1�[�P/� ���a2��ۗz��5�����0,c4��n�'���ߔ�1#$�׈�,�����z-ёes���:/Y�/���	6�a������N���H;7��!��]�<n�]JT��]�F�0��\ɟ-|��T�8'm�l��Ũ$����Ko�^�?'Ue<��$�J��S'�i��y���@Q#�'���/�K%$�����>Q��s������ev�X=���M��J����M9e�Ew� R�v[C@l�ֻ����hU���@ ���~>��b��V�oF��1���#*��`Eu�W$�f�.|�埆3pK�-}���"W�	�c˝��V\�Gad�:c�0�ZZr����u�*/��EPϋ'��E4��JՊ�G���i"^L�W5��i�:�{���l��H~��Πv"8e����ꥇ> �[)�>T4uL��+>M|�!��Ցd�)�󥗦�S�TK����=Z���~����[�?���uy��R�?W���7���K9~��|�OQ�R���JV|�m7;Jĥ(4�S,&~��tD�g�І��7ʕ#�y�zV�]/��� Ue��1��Cz�G�B�9�r7�9�_�Fx<��s��3�,����S���������RŤ*�`UuI�
�R������"�g�h�{�*$�w��z�e���N^�M8���� �F�Pa7a�$��l?��k�ax
� �@����=R�����ER�K05&W�Ɩ�9/Et�<���#�F�`� h�2jS '7!|�^ЮR�@���>a�Һ��"7n�qp��=��\��'�_Ԝ��#s��@\�,`C��mMo�T��U�ڻM�qn�k�ڠ��>����ã��UكӨ���sS\���_��Rcv.ܴ�\�� ��rG �vmT�r ʔ6<�����+�eb��ٔΟ�U���>�t�#�Q��e�Y����S-��B�z)ˈ��bA�Zm�
Ka{7!�UL����o�u�	H��ɘ����G�����V�W+��\��rѳg��	KM6��켬%�� �D�	4D����Z�@��^�����A��L"dt�bM��g����q[�Af���(јç_l�)"v��!}��,���ף�1��sz�[��k���e�VU�ā<-<U������ =C�T ��~{�:'b0F��k��P�ʖ`�)�*_�~�ݳ�)g ���$C%�=_�o��Q����"���	��1g'd�|��;6��_"�K�������P��h���4C虛�[�`I����r�$��`x��������9
�d;"�y|�QOͤQ(#�lͥ9j������S����}��%E��&�#W�"�1��ص����x�wYi�c`Ց��I��َU�с5���Qf�AG�a���cE�l�8��m���U��h�h���Y��bxJ=s��C{ ���Lj��s�����p+��џ29-�o�-��ؕ�;�l�5�Q��@ẛ��<{ZZ��il�jᗬFW %T�l6�P�?�	�Hpq����u�n �,C�Sc�/%�Xַ��.1�#
��Z���f���m/����x�pW	۽���5*|Yؒ�qK+�@��O*��j��F!����|�hm���uJG���g�
/�U$U�W����I���DJ��c����r����H�gG!Lb��/�G@���_�?�'�%$U�U5��渚�N(E�zu�����`��ow\��j��V�\@Q���&�!y�����&u(t���xѶ}�maS��L��;Q�.!��kzZ�T���j�Hh�Z*n����h���d�t�p��[���@{1�w��n&�`ay�5�ث��M4���CId�x`P6��/p���u�=��K�+�g�W����i���j2��bg����;Z9�&�����v�?�ɖv���y�a���� o�v���{c�F���m�?M�{���{����kC�}�Oy[���fi���H��$��i&ʯ{�o������+O�@�K^]a�L�,�skE���A����Ut�\�{M>:��?#tͺCW,ZO���AV@�4��u��]M��6��@�')��q�N?�`�l�"W��mO���)��Z��3iT���9+�S�޼�4D�O�U���P �y�q>���Б��~��EB�'�m�p>�3>N�iP@�{+@*�\K3�	��&e@W�:7Z}�ɯDt�Į$��ð�
E�`�Eb4W���=b��+�Gzծbډ�	�WB'��m�H5�>��C�'Ȱ �LZ��F�j�&����*�S�mӪƷ%r���y���O������rgM���̽3gY��;JmO�ķXOm��K;!|��{<� ��F�m߸-�*^��?��n�j/��Jכ�BL�' ��&�J��ȏM+� 1В���Т���i<�v�˲���1[�v>�t�:��k�8����c_�`���2�
�j��K�5�4���5��tQ���Vc݇�/@]��lϒ%�HC�y���&�ZZ]�=k�}}�jL���b�^傌�F�M��b��V�9�a�4�2M��!�%-ݎm����VQ�Z�,-E@��:��gd�UNC���im��V�����M��J�������y	�dM�L�aX�돨������hN���1���IP��!���1����o�e��I��?�0��ua1�Q��SxqP�I�P8�L{Bm�P�:�ʭ1��NƩt�ƪn�b�N�;�O{����p�K6���HA���dA��S�3\z����,,ko�G����mFv7�(����i&Kk�����0"!�6Yy��hg�AR(:_/���xf|(_3Xq������p�w$}��P����/�N;F犧�4��*�ZpP�q�W�%�N�4)!c�jѱ���n��>�Z�LSaF,�/��&x����Ʋ�Be&
���uHڔ�;��9�,J���ӂt����rO:#`YS���.i��о��L9JP�T?��b،�����9��������	C��ˑ�HfP&m�|��-7|b/9�ہ���ۮ�[2���4��7O���d�j�,<`9�D�#��iXݑou[�(߼�+���e�s��6�����q�㝧Q�B���Dނ߰����a�gк?�{_B�G��"����p�؇������-X�5�1�J	M0�פ�����fg�/0��?<Uo���`n�	rNI��� 	�!����&�����{麏�Z4��	�nB�!F��yjI��2�uR�n����Փ3(W`�f����n����� �� ���j�O��Ncxޞ��CT	���t�CP��yTZ�)�+�����@	H�k��6Eܞ����$�xK�b�Dm5�R
���݈'��Uo�s�G]&`H(̇f\KSz�Cyᬏe���
���K�sv��+�X�@�͙t��6�0H�V$w�M��/PL3<��vd|����U�~�A�ec�'�h����I�|2����SF���װR+np9H?o�;Z��`wP�����)qY2b����%�v@�xn3�\�����%�������J��H�+�a�G�_�WH3
��l�<���`Z�A��c3�C�e�;�E�����^P�F��L��4(Z	�f3��6��W'�Z=&e�`��Z�����à�|�Ԓ�r�X%�e�`N9Tw�B	��� m�Ѿ�� ��N���44����{�2�����KÝ��8�d��,�{g 볙�N-r�BK�we�&�1uh�]l�d�pǸ K�I��a��[�P�#Ck�,R�3U���ȶ@��pE���m���Jm�ť|�ݖ��kZ�zh:fCe�B��f+��Z��,O��ݘ��a=c_�0&�AT���G؉�q�j��� ��-���:6M�/�.�GF����)(�c[�$R;�,�ϩ�[�i�iHV�P�I���nKHٮHM;��J�����Q#��%-Kg�{��+���C�U��0l�h~��*Ńa+�F�8�Se=�2	^a�S�G$SN�-t3e� U�`��*�����p}=�0t&�-�e�l�����$����ck��p�r^,�S��К��ϭ~��4�3��6�����"c���	Vw����F�SA�ʹ�ꑕ��T�_�H<%ƨ7M�m�2XO�q/��&�e�?��,��"H�c�,m�m�M$.PW�[�>1�J���z��o�����W�US5i/�5�C�{S �C�@��Д������:w�3]T�6�D@��J1�9	�V�q��u=m�S\J���"շ%=ڈ��]�l8U9l�(䥮�E*�}P /�@���->������N?��-�]3ojM&� C�ѫ��;�&K��t�����p1��Gr��%����\�M�aXU1����W}P�W5qc͢���1I��)fi��Ѐl؟���}��u�J� =K \&Ԭ��8��Vu����6�D����� ��n~q�����<��HR�(�5 v��E��Ѻ�l��/F����}Z��a��Hr�RO�s�Q��{〒K�0�0<���%ߡ-C,R�l ����Y����Ed�D��.�4m4�;�j��/q-�+�m1�ˁ�:�j����T�sB�Xm��\�;]���2IWڝ<Lx����偄dZ�'�I�R%�;e�~Ll��H��߾b�弆_��C�,�6r�ōԒ��O�n�9��@5ϝ���.*z �����Wx���ȱE�9_kD�tDOn)V&�-�_A�ۻ�(��Y���@�4L�Y��-t�H.�3�J�����t�ݢ�(���+����uP߄�JT�Ĭ�(�n�xk=�릕T��SIoN�|�6H0�w�	 K�����Y{���'B��5ֿo��>���7�^}唼惲�,��D�}��l͢�-:��c�wu�<��'�E�C���6�����Cd"�싟3��*�8{��2��-W�v�UCބ�v�Ba�����MV�����V�F�'��XD<?~�lR�^Þ�l�z���&�X�I�^�-9�(���* ��f�HVu����Q��v�R��R�����M#��4j��9slW���+J�D�S��1�%��%���\CO�Y��O�?�R/��|���"�f4,�)/M�
IV��glN.�B~@�+����4an,��� O��b7B�R��0��M0n�QE��
pV����!�V���\�B��ؖI@)U��x��s�:��i/_Tx��/����)͜X�����*BWz��g����{��G:_$nݶT�N5���6�?�one��q�W�㥥#B�'j}�4�����$5��y'd���)S�,/"��8���D���X7x�N|���O���G�
�S�dK���^�+	��[<�DU�fؓ���6���'.+?#oK����a,u����֟���X�*~��T�9�,]����Ή~��8��ߑ�>![ڃ?#jHa�)��eq.��{;x�)�uA$e:48H�m�����ͽ9ɰk��*�#ύ��ba��
?Z��#����U퉯��"|u�@�ح$����̀� �G_�c0(�lA�ڐ[h���y T������OD!!��E�$� 7X̳�N��M�֟�n-f��T�D_����I"����6e��AE=��'H�%w���g����vю�����^�Qt�
�Qns�X�HcH&O_S/�4cw(��R��l�ղ�؏^�
��r��Ȟ��]g��ћU�I�MH0�����e��N�6V}�bru"�<Ӄ�q	ߌ!ĥf�N0n����t�LV���г�lo�/���a�nY����q��XLy���HA;�@LXJ8�)���$�Mޠ^��<$�A����r1���[�_.vN���Q����d�C����b�]��Ysg,v=��y��� X,�V!�k�X;��9Ԍ�k�r~N[R���l��L���k�3H�TVD��(a}���1p@��<t�奤���c�a'��[�����-v>W`�b�����O/�Fh��C(̺�5��ľ�ˠN��:�;_��!MZ��8�C2��M;J�����>>�=�'�$f�&ݸ�R��mZ $�p�\�ٹ�4&T�6�6�����$&O9ty`��'�i�t3=I���B~����1��%����s@r�n'��̚���5�B7�u�W��1]ۛ�WC馡τ�:�~_��љ�9�u�@4�a�/wrv�=��L��	�ѐ�N�=7�ރE�z.�Ů��@�4y�z_��:��&� ���� �5-�"(�
͑�u9ʀ��H��]BR8p�=_���xLvT���ЂG����p��0J�:��IIn��a6m+���;�ZR�R��5��!�.3�:����gΉ�7�g l(�\��a���F��M-�?��uK����&�
�<`I��D6wM��j!�����O�*�q��q����?�'C�����{�(����i)�p�ױQ\t+��V2'g�U�f�x�lN��*zF(�ߌ)�WQ��,˓���>gL����?,(��G�e(	D��}�V�n͜��p��9J����w���>�{�A6�[�K����<HA��S�!�C.Һn��Qe��3 .=߯
�)��.��5 �������h�E�k��`)��y�C���e�s��hσ�G�r��O����襡y���|�* 8O�0y�g�"�L��+
)���7z�8�K��`�fOj�N��;%���O m�̺"�Ĳ�Ú���&�ج�"�Eu<�α�of=����R}5:s%�#3IK}vj_U=R q�/
��~��o��l,o����(�l�I�P�JM���,?�X������K.@E������d��L�&�M�&�2���Ϫ���M�R<c݈��r�3�	G�$�fƱ>��q3Y+Ђ�֩����7��!��^���pNɕ�H{��D�Yl;���/}�&�bh��
S��*�mcrR�������@B?��v�����Xp�^� �6nD��&xƸ�X�����G]���Zl^͢ޫ��b� k*9����f����zE㧞�c�>�_����N�
�'ɇg&��5�
c�G�K��U@�}^��_S���l�����U��9D���F�F-}�eX�JB��7�L����i�y�nJ�3j,�)��ĥ�h3������/�寤���|�+�����<���D������W~"�y��4˳�����z*���XTm l^U���ʶͬ�N�%���a�O��_�� xb�G�[*�@_V�+	sn�s$-��
fN��B1<�g���;)4��������6�eI�oo��[�����cgd@T�jh0�ͷN�	�e��^G���d��4��h��^k��Zg����Z�S/<�AYDiw���
��bǰ���=+��5�^K��-�zu��Y7��EO��sZ�9 
A�1n�b����G��Z�����Y��?V�W��k����vG������"���g��,\]���]���y(ی�b�[�zF"T��Iܘ�:!��B1C�^�.�ۘ�[w0���h�p���5d�Ƙ�t�ٕF��=Tr���o3���+F{���0s�����T�S�2;
�_���V;p��$�=�U.�n7��'��)P�j�K�ȋ���&��n���R�r!F�r�f��Lk�F�� �}Vߥ#L�֒�܃�|�#-�}t��Y	u͛A��ޅc��
{GzP�"�~� �.����lMc�R�c2Y�BNf���"�����ˊ@� 1�C��&��s�-������]�FȬ���5B-�o>pŅ����C��(����{s+�83��}h��1Xƣ�Օa�tE"U��eH20Q�.�JU�%	��*�QV��Un��7�C ه(y,�µ� H,�5��@Z`�����B�A`�+�vӢ�^�Hc�<�֐�红�=�YN�^W��=0%�U�nS�3!X��q�db_�f���g=�c��e)Q�6�l0#dv����x>�o�:V��Mz���xq���_F� �[z��$��M�N�28�z�/z�j>35������rvlo��)f9���3������\��ʣ�.m�Ļ>cot��幒�u���G��d�R͞H���jʌ�p"r����["-�!�B�K{�֜�X�9��U>�P�Or��C	&���ȠS+��5a���,�,B�����:&���Y�����l*��j%����IVr*�t�{0������
�����Bcު[��>-%T�`�Ln�����ڒ����JС\��sߺ�\����T��q��M�wEpn�6(�͗��6%hU��S-lu�ҎbVx�Ej↛<��>�L��SU�/q#���`
F�
�Wν�� � �g�Ĭt��c��@9څ;������))�qb�T��c	�qx��Q�!�j5��i����k�ǩ&r�;��"}S�%�Vc��R-;��k��*��-˧�� &'��x�N����2W��;�{7Ob����$�9�>����N���Jv0�Kj�|�7�l�t��m���٧��a�|���12V.�g���ɰ�0�F���T�A�;	�����߮�R4%�`�GJ�㼳P9��9��T��f����E*І���-l)���9��%���� ��ް%{~����9�m�	y�$Έ��ą�#I���
�IN"���c�ta,�l9"G���<��>Q��5nu����ZYav�+^����;�zӰ�ln��P���d�x��b��&��ˑ�!�U�?#\_�3�u�_�+X	o]d��E�M���B������p����goA����MR��S�u�R���ds=%;3�[�Vncd���24K��d�s+PIi�H(N��s'M#pUXI@�F�:F��Օ�_mL�Y�q�S�:E�"��hi����;�M~;})

Q|D�L�q�Ĕ�>!��bc&n!Y��*6�����I��Ez�T.2��&��f��_�+q���\����OV>%�;Od�%�&�"EL�fC��f��!�?��զ�"ԅG'g~���h0d�3�����zI--�S�EbҲW�I[��e��T����2�ɛ�����uB���
��F����Cu����i��B�O�|U�r���8}���lLo�Y��MN��H�vI={	���E�T��Q93i�ni,#���|-�/��1=Y��Gּ�sW��x�u��ULVh��O�]�S� }E�A�aT��܈h�Hz�]*�_��?G�\aFz��硾om��ܿ�����"���X,�}Z�����<���HX,�k�H�����$���$�T�Ov�ش6.�!�Z7#%.)�@&$ �>����J�G�-X�4��1&uS�o�����~��L���~s��n�٠͟�H��d�O����R�:/��r�-��ڞ.����{)����(���'	AAC�+�B��i!����fxz>M��ߏ;"��#�� �-*>T`_�8�t�2g%�Q��gԮ��w`�|�zG��p�\	/��Gː��_�HL��~����n�Tk9_�5?B��/�$�*��u�Y����5�.13
��#�u�2T^��ண2s�Ɏcj�.��v?�E�m�D'=DY&6"�����{����44��@WO[J��Җ�ܺ���b^z��c�G��M������d��t%`D֬�<�7�?Gf�nI|�A�+!t@���d62�v��	���Sx�Z?��	�㛏�9�s��_�����lT�"���Ìj���L��<� H�~a�"9�xe�)C�N;��%ȃUP��	���C�\����ͭGx�X�Q�#!�)�ʫ�lqjVF��ќ��,[1 eAmU���v.���;L�%�dY#+n9�������XN��lZA/�?���T�����k�:��Y�t��WR�$��U���reP�֮�x�� `������7n�Vቐ̯��Yy4_����pv�������"[��]r�>0��-��].����R�1����Y�0�A�_���.C�yB`�G	�U\�i��.xA��X&@�7��Z�S]�V��N��W��:�r��(~�FaU-ۈwf�/U X�ѐ�%���Xvo�y?��Ƅ��z�;�_|��k�T��$�m���U�9��*TY���UF��ZM:-'�z���kX���j9�k/��ֲAg�P\�x�.k�u�U#b��(�U4*'��C�} Ik�=@ǆ"~]k������,�!�����E�5�JR��h�KJ�����?ŕA�ꪟe��Z6k3���-W���<s��
����8:���Ώ��<��	4u��nBp�� ��t:��Z�1y3�RG|�րy��=iYxm	<� ���j�ҊT�y��U�t�yZq����\���U���FU㋀�V�:R�Rmt�0Y��&�ziLy5s�D�;CO����U��5-�nZ�3X����-���� ���b��L٠U�������|\U�q��7��|	a�5��X1Ĕ�ˠ#�)p����Z�ыS���ޑPVk���:�4s�(a*�S��=��V���
F��;I=uL�X�aҞ|dJ��=�M���oO��ڛ6����lž�f?��C�߫�}ۨs��U&�5+����FI����{���}VD��u���ۃu@�(4@��Vp��y�Q��RA�%K\��t�;pQR�	�i�1D�3�cY����`���]�қ���lO�3��G��٩Kd���S�otՎ5��jΰ��5�f븐-[hފ&X`����	�����E4~�$3��%�@(�ڰaP#��C1��Z�^�?�׍F��kZ�jK��nlPdUf+�ot�s�E65{��'�e1М�]�%n�+��¢��#}��m�c4���S���ɛ�Ǡkޖ��)�7�0���Ų�<)��w�(�?�j�Õ&��-�����u�5u��T��1���ge��p�@��Xu%�l�zѣVz��9���ęʇ�/=@Ɨ����َy��:�<�&����p!��i���]�R��+�V�|F*h*�8���+i�<K	/�t�φ2����_'%���	���A�J��I��4!)��RVw?ruq
Icd��#Ѕޛ�� ��_n��&%U�-}�r���-r~1��K���T��S85ҿ�f.@�����tJ�����
"g_�m[�c��WM4��]�i�c�7�Z���]Pxk�zt��^��2��|��]I ,Y��]x����֭Q��)�JF�s��;���ns=1]b}���
��dwh����r��	6l���3Ke	..������o*��le��"�<R�P�ȷ�=�����C���F�E_n�ܩXɋ32[�[{#n�0�@�j�U�y��\��GT��&��+��-���ɣiÝN��������qϐ�b�+���1��>�>^�?�X:i�ѣͳ���/aN���I��Q~�߼���@Q�j@�:��[�K�lO�.����c�w8���0;.NZ��s^~-O}_~ϡ�Z!ۂO�.-����Ǌ�6S�����3t��p�[g��䨧kl�N߰�`�z�'o���i�	�����)x�?��h3g#D&��duY��VqG9A:����M"��K��"�8�I��ܙ߭�D(l0��A����h��P���/�8�q�<C��=EJ˼��d�`V{����beεk�Ζ_��%��\�j��e���'�)�US�R�ȅ� I����
)W�V	Ks�ֹ.K�^x<$���芡_:�n)�ʨ8������+v�4�e������}�>"�mpN6����S�0���r3v��f�S���:��3��Y��&hپrP�r��r"�D)pPx���V0���+@�I0\��LF*3[n=3s&��V��&~��o�oH��2��~}��yt��Z�Ġ��p�-�U��+��7��&;�1��m��~~dc߇�g,/���g�s�*�̘�
�o�/��'���ۋY�Y��D�7	�<%ӂ���������_m=]�Jw�%BC>W��sdj1�$��(����-�`��:��j��P�!b���v��{-��ˣ�ID�n���i���0����F�B�?��?^�?�����0�Nt{&d�u��r�?蓌f���wB��F�]mv�f�

R,!77��A�Ȩ�]�a5��ɾ�;��F�\������2�j��\��x��)�L����}��NO���������}Jҥ�iJ�;�č�#�:'�C��z��;8Ӓ𤋮�D�,΄�)���*��%KC�"��*�R��"���Ҏd0c{�
�9r�p~�^J���$����i_��#����z�ְ�f۝E}�L���>w��QX7V� Q�?�z�����\��9��{�w����Mk��|�B[��Wqfif�v����ڶ߼;XmJ��M!QF��۳��r��S��r�͎�Q� T�7����,��.X��Ǡ�kf�>UKq��[�V2�#�@Ή5��5�0e�8�&i���8kx��@�8����/�Rƪ��O�)���dk��|r�����J��,�C�G d �a��挧�B�a+�����N�$��+��5����%� ,B�>$-��6Y���`kD�H��$�˖L��;%ժY:��������s����w?Rg�5�;l�?7JTFL\˥�X@�j�3cv�v�k�	���n�0Yq>b�|LT�d�y������8�2�#t��1��dI�H�4х�T�z������:{H&���:��HG^ �mx����G��ҢdqԳȦ�9���d��G��:�v^j��<+�o`�W`Z�D��1�s]LG���e�s�Ǣ3���Ne�AZж^.�L)��)wz�-�V����r��˴������KIp�GhYќ�Y�5��E*����qQ����	�r��zAq�V�kǧ���8���x$CsC��1�kR�Aꆴ�m��XL%�#�����Ӟ/��c;���њD���̸vd�7QԸ����ٸ�5Q�Ya!���C	LUʠA?מh����a�ۓ�O��ꍍ�Ll,Kp%����|�۵K�*R{��M��.�I��:�������s뾹�_ �I�<^��<گRȅ�oAҰ7�nymn�'�hz���;�N$Q�U��V�)���3��v%���͉���p�2�
oZZ��4k:���9��.���'�Z�3��>ׂJq��Q�ě'/g�U��4�J]�g�W�;�����<��Dq]� d��ƪ!�.�4�No�u3w���k�=;�}}�ƕI�Y�]q��D�8x6��Жu?�S;`_��IP�G�*�G��fL������%�Y#T��)3lʅ�3�V-",�#�oi?4d�mO�w�+�տք��A@�u��	��%��]��-)Nd��.��LԋT&?/|W��3)���(�-+�"7����L�
��C�
^��W�;�&�^R����vJ��F+���V<����v�:!a.��qM%��)W<X��izE��7J�����l��� �n�:d�����1����NS��i�'ǻ2�o-f��P���|�l�)�C��	�d��(�X����i��IU���<
�*�����]"e�<Zܿ~}c��{��2���m���X��d>���t�_�ٶ�l��&�S;����cmK�j�Q�zۚ&���Ҝ�2���.~	�O��¶���p�bj��1,���]�8,��a�F1#�v�_���v[S�8R�D�]5B���l{/�7q�D�ɓ&�쫥4$�)�麢I�T�I�C�o��ΣO�j�{���}��=��¯��s�%^��J���b)ʀ���3`֔0���C�ɽ�n�¯������C�}��e��uO�'%�������W������HW���u��։�j�M���wW�(�>5�$J���>9H�џ�إ҂󾖭iq����@�r����J;��C����c�����|_Ca�g��U�'��k�V��l�Й�І��pۇ���%�/}���E`˱X�����eTL�뎊�����͡�B�()B��um
�;��O6��n�_a(T�lsHT� �Y���qPDc��(?,�tŊ-+E��8-��0�H`?L/Y��������J$���G�V��ve��㝓Gt%=iW(x��ۜ��L(�����;�A�v����&M!H:���h;O#�%�t���"L�H�����;�8P�96~�x�3y��\��������X$<�ة�Im%v
ԸÜ��ᳬ��x�v7�p��5����uЀ;��sEh\e��e���*r�ȗ1�{���V��������w$e����#<�{�@�
�Ƭv՘a�Xk=!\*Ʈϳ��65�����|�7����\�3�@���.@��9�x��N��̿pu#��Bp�BC�o,�ݚ�OǸ7�r3�� ���h�J^c���Mk��|�� `
��;+<2Ĥ������%�>�=E�#ykI��w�T2ݝ3=�e�i�r�c��_���y��k�yY��rE�2���u��,�o���eR�T4ݧ�lr�ԷI�$>��|�� \6YA��!��F��H�J���%!����֧b��E�1����e�>� ���{u&/��BЉ~|������P����0���� It%|�F4;�`��C��}vsB��)����Q�f��:��s���܎����'�'��9Z����!#ƫ.���w�E���m8�w���:�c�O�l2��e��o��)��FV� �S11L=�Qb����q��,����E !��-6Ĕ8�@_�v���q�UV��q�����]��<&���@MHE";�Wu.�4�����NW�l�?�h��A}�N^�u0v�Sgt>h�`��-Qq��F�"MM���3e��z��af������<��J��;)nYi�����>1�IS��}a��h��;��1�k���d�\��L&�dU�e���m ��Y���4��lBC����\��x9<5��dDo����1��b�8����k�e�EVxXJ��(:�s����=h�i5��ˑYo W���Ӈ	�+}<umocS*�p��jp��ͬ2o��$�aH? ƍ'����a��*c��z��y�'�lQ��m�8�����E�jO���#�*��}�7��q(��c���jȼ�C�A��J��6�Rz˛� �2Z� � �=KJ���P=�k����}��n�	NJ4�,���^t#Q]TR��Ÿ�]�B���g�w�`\ĝ��)f��śiZ��R��7���6 	�{j`Q�q�HY�-F�ʥm�#�v����1H�P��V8���ɓg�5�GQ�������.�F����Z<���Ҋ�!<�^y�p|�l��Dw �Y�|
,���
��Ԥ#�[_]��̎��E�3��HI�����P�fNȄl̉&M0��ǝLĕ�ع��_5G��Y��J��<FF��b5�Ւ������!m�J�ۘ�M>�,��K���	u���H�]	U�A���ӎ���N����38�O�T�;�̺	�B�p��ZT��x]P�B7O~A�}�x�7l�,�'M�'c�cE�����o��{�nJ�"q����8~_���q���BM=����w�5�N*�����3�p�T�F�h���. ���Uc�qU#kI�	)4�<�^N�;�:W�m�'��t\��{h�93]�O�,h�P��l���m��^�wW��	I�#t\���:��U�{��g��R{B\��j���s�DpkD�^C�Io ����`M��Q���ՑX�c&u�.�"Ma�����[jr�䨈���7S�6���L7c��nSP߶_�MSm�n�ˏ-��b����D˦�1���~Q�	� V9vm�dl�5>H�
8�s4@���Z��0�o5jz�.L�7r�A��(ذ�5v0�/�g�v�6$��nk�0�xn�>6A���@��M�E���,�tquzVz��~wsܭؓ�)�����.v}��SsU��ۛ`r��'a�ܷE�u�\����oO�"#�#���8���H���z�v ha����zf�����☩~"8������=`�\�_K�ǵ,��D�.y�[K~��d�]6-�
�Y�8���<H�,��W��W�FJ.��j�"@�v�A��U��a�i���_,U�箤�d%ȵER���)�X{"�%���gYUlW*���,.4,� ͇w[:-��R䚁��bZ_-]�N"�A�+��U�@-�d[��5��JJR���P�K4�ď���!ζ)k�|���F���"ƺ�_�|�;P���.�����xӲq�,�P���J���a�--���&���fj/�0}*R�_?����X��"Q�>�\�w�_Q��%������q��n���
�k�>��iME��חN�g-Y=�M��i��|f�3��%|7��O?
��\ϐ�B�!�fr�?���g34��u(�^�l!�uf���2��J".a/��.�((���,I eM����9j���:Гl��!X���jx�GR�ֈ3�c.ʲ�>�  ��o�lf�?E�Q��o�1��^��b�,�Y����AҨ�k���������2��V��O!�y,O98��R1��i۳�6z8m��Jp����$D��V�O��1��^'x2�$F�����S��9�|�A�Q��;�Q骥���1�>r%��IRi)Q�[��$3e�w0���qO�oOH�D��`@���� ����,��K28��Q����dO���a~ؿ"��,�;�泻�\�B��mWk�_��ŝ.r$W��3�>���T���ֵ_M1!J�]�k�w�ͩi��GJ�(�̀�#��zx
�y�� b���+)�0���W߅1���da���6��x@JT��:Z F��7
d��gϓE��~EM���.�bG����:!��p�/��Sh�
�d	y����0s4gp���|��w�.%���o.��O�i�n�K<���,�*ɛ!���������ص[��)��3��+CJ��"�\\B)�m�H�Agh)�V��Ŕ�]Izɞ�K̈Iv�5H�v�
�ij��)���sZ¯�c����I�,;��G��5a����1=N]:���gLj��d���u�͌Γ��CwsV��O�C��W��U�{��%�-(��qd+��#��jì��ȟ���㫓���������ϧ�蓪�~�fLM����?���ũ�s����g^	����G�Q 2_�3����|=s7/S ��	���>r�S�ZG(�d��a)#T�Eڈ�  Zꍹ9z򴉨WH���A�����8
�P�hQ"��c�dK w��5�t���g�	1d�s��ņE��7�_KU�*R�r�;�L�% �7(R�4��l�EC���woi�SBH~Ҩ����u��=��l����2���Z��ǋ�d����g�k%*=��}�+[pY���9WeJ����)�Ŝ���G��z�>*�|GO+(t�h�|}�4��lz����X��Sg�xm�}��"� �M<�rO�Ţ8"mZ�'ߤ�Ag�e�����������ȥ�Sr���p��⑁!H��v�	�HCjCd�T�
���S��'��x��qRFu����%��-��g�^K��V����>.H�U��#Sv��c�VFf�����td�k)��^��JH���%M�dD�L��D�DcgٶS��ף8݌$���H�F�mZ��g���z�X�q�By�*���1��%�2�ͷ}����Y�5i?HZ��_3|���z�Wn�(K��5���VA�+����a�;;0�d%��vI��~���Nk�хҁ4Dig{��G˶���>�Ev����c9 R^|yL�<�~�WW8�֞�&�Eb�z|����,N\���ƃ^l�^\�uy��j�W��>�w�X#�k@����߫u5,O���_Nu0�2�R��AK�s��yÊ���x�uW@Ohb#fe<V6ՙk! s�!:�B�m�U,��H2�|�w󪨓�8���6�� dTT���da��	��ʬ�0IU����bhO��%Ժ��U���h�B|@�Yr�T ��Zzl�c�w���ʶr2�Ei.��,5Uq?�A�tZ�H�s��-jQ��"�b�,Z��y�`>�Ι�P�F�t�k���n��0��A��2P8����![�|�J}��6^��j��H��6�fˢNVJȒ>�"a2��n�}Z���(���6�K:kJ�����H=߳(��j���?���RC�������"����Jh%��S�>\�����/PT�3ud�Uy��[��9�/?�-����츘��.�	af?�H���0p�?>N�x5���@J�G��`.+��/�E�;b���z�E%eP#^� ��ɓM]�e���w��no���V����*���q�M���<E%EJ̗s�lN�|�+\i��d�5�x/�8��Z��=�P��"'nX_j�T1�C��P6��aʃ��®�=��w�mJ]��.%S�ڈ��&0�\#O@kd0�v�
�d�����ܳ�=�\¾t�'B>�d��ؘ�R�A��edG�8���;)���k'�䝻���f} C�؞:�Ǥ1*����II+��m�1*t�*_ x}��D!�4�
�7��׍SoI��+%�	��<f�7UO=n6��'D��!_�kD������	�DJݤul�0���Xϣ�{��w�=h�b��x�w���ka�CI|�.��l\��Z�0L���Tw�+�9E�Dkж��5��ۓ���;���FRd>E�χ�u�6���c�X�71�(L��-+D�D�"+w�/n�t�>����!�S��$q�nlБ���{�Pq��ܸ3�7k0,{묥��h����푏�rw���1_X��.)����t]����G��Hm����ɝ���>��>Ay�î�%�r MF��T6�73)fHQ�xʲ�=g���:ِ�o�M�vI�$�����w��2��POј4�
������T�^�Z��9�	�ޡ4�Ó��4�W8�`!V�9'���,@wV�j���<��C4D�N(��5q�-�.��QP��\lLU�%�Z�"��`=�>6+��U�Tԥ���;γ�"Z��o(p�����C�Ҩ�G��_��-rצŮ��%�bíy��۵��c��.����0�r���Y��/I�x������R��;���=��\nFʈ��U�X�R�NLG"��Op��.MaA��uc�R���_"�擪=jA�{m���Dz����2J�z��Bf�Ce����J��p������<^c�M����_�ڥ�H�4��1��7k��L���'T4���,�q���p(�H���U�C���bx��b����?���[�R2v��@���)yF��>�s�050�4�����%��S��0{�g�<w�*mɣOV��A��r�����a�%26��v2EKr����Q�L�$�r��
e�MM	sw��K���1)�@0wx��6�B,i�{і��\oI�N��F!r�/�1��y]/s4H�z����\j�}OӚS� �j�.�*�"t���XL�K��k��
�\���Ľ��q��X��:���K�w��'�&�
���C	;8���>v��h�H���k�jF�[鼙k9W��A�*Ӏ��f4=:�a���_� ��N R0{
�����o�O6J���kW/�bD���0L��`��B��"�ZC��:;K>����/#�!w�U�i���j��g?:'�eQ,��� _���CVL�L��oY�.2�7��/�_�pw-�7�h�W��3pb�8��Z,N��u>o#G��$��NzYK�N�L�Z�����"��6)�oq3�%Ǐ���_I��n(��b�z�vn>��C;��([������k�:��_��~ח�OYi��a�����"	��q�q��W)%Z��
-nF�Y���g�����߅@Q�����y�� �o�mjF�7t���-� ��&�0�+�ݕH���K}��5��U����nWR)6Y��`~x��]�kYk�3�	rD�ڜ���*�.��顡U]R��EV1ON9��啇f)H &����Ei΀��·��;z-���+@�ńA���󰋳A+d}|h1����"����a;��X.��v�JO{C�z�2�|�u��i�,��"u�T�Jx�PC�=k�fbd��J�/��m@�V]�%�ڳ>��u?<�?�7}�3;pY��z��Yg�v�� ^$ٟ��C��Bd��@3����L�4����)S�N��ʷA��������>�w���1N6��͠AI%$u���D��U�g�#�;ێ��PC�s�Y3B����!�����^��d|��UQ8e;:���x�ѝ����0�����o.?�O�����?�@p���*^�3լ�7Wb8:AfJ�C��'G��)�~&�͎����DQO��:�"�7�>�G����WTj$�=7�b=9�$��/(o&N��><����Y%�o��sN�D�|X�Z��$����2K\���U�pm)�R*Z�أt1�f�l.-�N5&�jZb}R��5w���#׳@E����_C�¡꬛�Ņ0�(vr��u5 )�Pr9²&^��gK��Z��0�[WeK��a�]n�+�[ �щ>�-ϰ677�ѫ�?�����)�bQv��a��9������;�j y���1���<u[�=76�R y3A��K��Ә�Fm�h���N�t{O7�F��m�v<d���n�X�Kߺ�y:	�+Ėi�D�@�;���1�?�]���JJ�����HQ����~�;;�F�\M�xP��4���*�l��i�l��P�&�_�g]�7�QZ�FŐ[G�e\D#�zĲ��r_ +y���%�:��R}���u�i�Z]��d����O��m��O���2�[�ڽPk\���W��Hv5�c���󶏿����*N�`�Z��848"��X�9��M��Z�������,�ڂ����t�D�L� �aX&����Lr@�w��K�T*�4..��ߡ��8ֳXs�4�B��V�ȠO��b�L��I���?����zz]]���saUW$�ÿ������v��S5G��j�S��)/��gAI��/L������I�|K���#�������=�O�����M�sD��7_��[��A �I!��`�R��/<���_���t�d6�PA>o#L`e	!��m�P�C떚�.mE���e�qS� d��g����+�#�(%'��?jv/��&�F�=&~��A�'�3�r���K��c򥖏w
��i��W��Ћ��!Y54<*��U�xjFf&���{T��sN�C)���xř�m���	S�Q.�k�u�$W�;F@ćXhI~�^`�������]�QC����_Yc���;�Z��3�ev�_�z�񎓝�n�D+��z�P���Ȳn\�k�*�S=��o�c&v���dd]�d��L��d���4�YC�3O�{8���Ȉ��G���#�t(>�]���_�P��k+�&�;���:��ѻ��!��<�����T�|�����iLՙ��H��5ጥw_m90�6������[M�\w�x}s?��%�Q���C�m��� ?dܥ��5\ԕ��i���8Ɨ����[KqV��#��"EqJC�K	����i��乙k�+�9z������f�����"�bs�����s(�.�z2\㦥�%�?�ӻ�e����a�pm�)�Ƚ
Xe��]��b�~�@��׊�sa*�}�e%��8�Y��#��Ʈ�s����1�o��g�]���9�<ߧ�|�:���Qс
W"�����Q�;C׺2�!�&��S����[n#$��&�(�$>r�	d�ڦ�4��aې�2�'B�튫�CV����)D�����U��C�Z|���A;��C�?����U��l���e��{t���!��tj���'�Eo@ub�#��O1����]s�7��=ݺƣ�"?5�����,OE(��ʆ5cT�*�Q�v���Tw��L�Ԋ�*���� ��] Jpw-�gP�.2�x�o�ix�h�$���ݛ�f���f���IJzA�.���)�8"/o)��G��
!~^��M��?by�nE�x(��l��2�<%o8;U��U*UP�[��篢Y
�B~yܵ8�@/Z  E�f������U�-F���R�4�`B�����h�Rv��#�ET \�z����q_���Ƅ�	k%N��ƻ#�0��?mO0�����,���48�qWw3�����!���1��"���J*!^�Ϩ�&]ܱaRV�4�e�n���sm�"�!C�y8y�=v|�Ȥ5����*�kY��OS����v�H/qS���i��z_W��O�7��U5��N�O$���H��|��#�$��:O�$�KW��nL &�v��'�3����Ӳ��)�F��MFǓ�hE}��V��&f��c���GQH����C~8�;�M��e������q��MwK5O�1_����W�Z$w�k=u�p�ȶ�R�G��h��sh�X&���}M��Ni�%���*+�*�k�z>]� �Kϣ�=/��s%>`ɮ�`�nf���b4�dc�p�qό/&��(���Y�b�Ow��'#z}���������:������=����δ	v���ca����LJ�Y~���z?��Է),���.q}�\���H��I�]� fJ.�x��!x��3h����s1�B s�g�nv��(�I��0O���&���F�[���Ɋ?#|!�ig���*=�Ԛϝ�9�����6�^��Q
'���y}�B�����»��6�Y"��Y�N)�B���&�d�)��W����,������b͠��UL��ʐJ�ͦ���&����e�=%���Q 1���e�?-�(!�Ny�t�w�,����`aZ5��5��9��Z~f��&JTF��+Q�㠥q���y��V=�[m��cS����@��f��P,��^�o��"�^�u��fS��K� ���#�Ln#?���e��4j6Z���$�ˌ��ʹ�a��j��q�q��K��,�Jan���"����[�?�'k�Yv��×v�ɞV�w`�p_x���\��y5r�����	�e�z#�LRYi���z���C�beJ*�Fpq���=�`�!�D/��^;��tЎ,pZ��M>�,
�8A+��ו5��:R��p�����~�z�`�so�y�bM��`g
�D�@=���2E,��l�D�C���?*!ӛ��@�ߟ���(��K�@��!�Νt��e�RV��-�_�#��py���v9vRY�]��os�|���E`���qa��y�6�'���5pJ�#�1�	��
��/������1�7��q�����L��[��o�H��!�RS#�u�]����D��؍�?W�����p7;��P�Qx���th�k)~����D���V�d��Xwsk�y����	^�e�ۙ��]������(�l�U�/6m�J(���:x��ՕХx@�F	�e��2��Ԛ /6U������{i�/���4D;���+�&���7;�qe*+I�2�3>ъ��@� �Ld}E�
�c�Z�#I����}O�+?�3�D)��
l8i*�e
�9���'!�����η������6ON�{q:�e��R�qJ_S���%?��c������{�39�O �F0��M��=�<�������%�ډ��{���KN�y+��@~�2��7,�+�s��FE'^",!���U1��3xκ��GcC�J$���v�v��6�Ч2���S�*�-J�?|�5"γ"��S�
E@���~����.j�H7q�@��Q~n�����,�E��L�V�uëF�3Ö�Θ�p'�G�IX}V�<U%����Yی$_�MN?��70^?0�ӆ.� Y%�iK�����Դ�������D�a�@��};�I\����n�Ϻ�|ş���I�����#��W���r��|���35�|�T�"׳��|�{C�f)-��&b	��:�!@:�n��ޝ�[�1f��n?к���ݜ�(`���b@�gQDMBJe�$�c��u�vI�E���+ܧ -1��v^5�Jݩ��Y�a8��ϸ���R���'y$�q�;�n�{���0�E���T�o�V�S�LY~_��2������htT�xe�l?Qw����o�q�4� ��X��o,�MIv`�4%�-a�m>{D�6񛤆h�r�־��x����9[�q���8���ls]e/��o�I��,�t�I�ӀI�..�	��	��)>=�x�i/�
`VB��~��
Ұ+y�"�-9[<Ϛi�ƒ@y�a�h�_(Œ�)Z��J���U9�3���N�K�jce��e
~#���hw�<����¬'�)��C&�b[hqc[ӭ���[�����}���DG��Pa@��F��Ma�7��� ���L��q��z�m�"?N�a�E�oq>E��/;�Y��Rx�e��kf�,>`="���	�\d��0�z��dXz������5�~�`��ߐ��D /�������٥1Ђ�_���(�,��P�G����$���g��e�R��L�z�S�[��Q��'WJ˪��/qķ�z����s����i����ڻ�]����N3s���[��0���,����h��z+:5���N~&.S����	�ƶ8l<A.	�'(B���w���=h���� ��xi�1�q4�X q��yi1�����L�)��AQ~�����Mzt����y��.�����d�%h'�i|ev�Ɖ�`.֝�O�U���E7���]��#a�֕EDP��K�]�&�,�\c��/3�� Mlu<�z��jK����c�ޑ�[��n�4��#/'��;Q���g�	���l+��?�������owHj�V��w���0�L�E�j��60G�*������t�5O��O؝��+�<u���ْ=��!��� �uЊ�"pGA�x.����;��v�x�8.�[�Z ��eY��v��4���{����f���ݖ�D5��ć21<��o^ℍ�Ç6�q^�Qc�E���ǉ{��~���=�sϯ�Ͼw���q�����8R4����?e�*I�kbM�R1�#.Ŝ)S��.Em���uLY�||��%Kk��9ѯ	{�i:]��Iv��(f��b�G��&#�%K�}WJl��o�"����!ApIx�T��/�)�n'���|JW�6P�:c�-DE�/DT&�U%÷�+�8H��sv9﫣�p�u���Ԅ'nܥɠ:�)�ZEM|��"gK�v/��#���8%g���߄��#�"��ZQ'�PE-!1Y$pW�M��D~3�M��͠"F���w)Ӡ�UT�U�[Cr�P*mA�ԕH���1Ƴk���i	�V��Pm�;sZ�A��46��,�m�il0�sm� �]N�H�/$t5���2Q�<<Jr�Ƈ��W=��S�/,�4Y_' M$^�O3\�
��Y<pfKm�W�&H��o������!	��0����\�X�礢�1�Eߠ��1 H�����`�Y�]���`�-�� ���1ΐ�O�hL��N��*�k���U�@ٯ�KQ�n[��d@�a���k��>_�De2]��M���a\6��/"�h����LmF@DH�z���uE8S��Ls>��2h�L�s&"��Ei3��8�Ԭ��Ro�ߞ��F���hDG�f�k81>Y���@Rʹi»#��a� \���F���F5@1a��◮�E��Adr> F{�+��yG�����)��̓����]�U(�Rit:��Ix�n�@jd�.�m��>�D�)��/:�8��;����ڏZ�y%GՍ�,gI=Iw�m��=��u�RVܐ���.�(I�%�Uvk�fO㉲Kٷ6;�	b�[}�]el����>��������C�lP���f����dAR�
�(����^�'��.�灾)j�V�ULĊV-�\�Q�'��"����S�B?!06��(�����|�k^�^�s�R���>��Z�]��N�a\d���P\8h:�ƀ�0�-^L��QW�3��Q�RQǿ���g<s]����Cc��	�}_�-x�xy�?>ש�+{>�I���֋k�[�j�˅�Ĝ��C>��� ��R��=�	��s�G,�@ܐ�1y*vès?g���7�ZePK���M�
��`R�C��<e�VŠ�+0�{C=���ӗ,V���0MpO�=={�݁6Jr�^L������Ĩ��*�8�^G+��5��%%�K#�� ���S0�2�Ц�-�шk�J����Z�i/ 
o������.?k]����wU�IH�c�x���@���î&�?vV���\*3a������vB�t#�;VgK��q��ݾ.��ɸ*��&+ӓ���@G����An��̱4fXd�5��(oN�O�1ye��X�k5e�j.�a�n!&Rӛ�����J`(r]|aK�K�ў^q�P���� ��/��^G�����Rػ=B���M����Zm��.U�(n������Mr��jA��F�r	�2�LD�,�w��L,<���3���Vs7�f��b�ţ]�'��V"��#�,�*ٜ�n�V�r8K8iE�x\��u!��k5p�|K �$��2T���r���{5�[-ړ�P^�@_�tD,��X�];�$W\�")HI�ژ:3Ds�>��h��K��Kt>l
='��o���u��¸���3B���o��JY��
M��%���b��y �L�(%VC�Gd].͠�2 ,>�h�l}Fd���X�h')	{�D�p7��%�U�%X����V�ۘ��� ��P�ˢ���ʫ��E4��P��3����ӕ����;�3��qǍ/�T*�^�]Y��0Ӝ�a�j�vfm��jX�xy]<�
�w��*󮛻���|nH��&;&� ��ct|	�VT܉*M&��i{�؈�SE��R��!-�qS�"��¨q�p��ur��P�`Q+����҄h¸��Z�!�����˹ڔX��V��XȜ�TIڹ�d������l�ϡ�:)�^�|�����²]���Ȥ�j���o�8��d�v}���nM���%��*���8�,�Y련���%��:��Z��m�ˇf�w���U�Az@I��� ��~����!�'�e99�}t��I�Bl�9�@����v�t����kJL*���"(��y�D�}�%~N
�CD����t5D�Y�u�,�dTc�1��\.��i�`s\����k �~$5O�8[��Ji>��lVͰ�4oEM[z�DW८B_�CبT�=B�i�I�V�Lco��&u�R�A�>�a�zI�q7�/��E7�����1���Xv�O,�Ipoe%���%�n��K��:�&���!�?�~s����vx��VV� ��jL��F���nO��I�kw����&�H� UHT�*�rBAO�]��t�J��7��\�{�3>r���f�����H����4ԂJ;W�~\]�wa�t.\j+#���JPg�d�#��2�3 ��7����1Y��ѽ�Z����s�J �p�vԃ�� b��a2�L�~c�s��>�y~Vѿf�ݠ�"O�>A:e��q)��<E�	�"��N��ם��}�� ���\M��o�Q���K8y�v㵟a��)�ƈ��wL��G�^(��?qTѧ96M`��뀧�/��l��i
4&3�K�g�[ݧ���+��xE�QM
t7}����O�f*����qf,�����@@�{ꊪ;�Q�GE���C�G8^6\+����5[��rds�)�Pk9��k�v�A?V�=K�I����o���^���T�Z4Q�I�Esʭ`�7Q[�����/汃�@�a�sf���$F�^�8���NO�+�O^���K�ZEbc|�!�T*+v/D�̒�T�pwb7�uz�<�qpʆST<H�UYK�e^EZ�etwA t��_�S��9x`:��`>��ɞ`�ScP�&r�k�0l5�|�Qy����J���.�ɁD��i�ѠK����a,tl��#�M4+@)�?�1��3��
<M�=��eϹ"�Z��/���2a�.�T˓[h�X���� �=�R�\����G}�n��������ߝ��0wg��#1�Gtu
Tr*�Du��M~�2����6���|#Ƞ몀k�������60`1ҥS��W���:#c����� k[n3��)���b�wX�OB*���6񚯂4�cz� �
1�{��e�o��:��x��!VʜQH+����&������c�U��{�q\C4�E�*=�B`2��Xb��͛B�� ��W�x�8��A�#a|�ζV��V����W=?^Tr�>y�2#|��ko��q�Y��5D��Ӣ�5Ǒ�>�B�0^
� Tc�i@ۛԤ llP�o���'<3�vŎ�|_�o�'��{�K<��(�3q[�a�5����gW�K�r@K�����i!��:)D��V�c�|[.#L��X�|��6go��ϙ��z�����q��>w� ��0S�_X�Ի��%� [�*�%gΫ����v=#�=�MRi�O��	�'&�̒O�f1��[%{�V-�Z
�k��:wbn��J����da�4�^�h\� u�V�,7�h��#7�ѥӄ��Z?<�.�#;�K�(�K��K,�C�8��2�9�]�U� ���@B �V��&1�)`8����U�$�-��P���X���m��.I�g�j�	W/�y���)|7��aP>��S����e%tog��Sk�ؕ��a�ݨ�	��2�V�Hu8���T�m�q
+�_+j 
�N��,� l���8�g5k
�6�7�̾�����s��]�O"`B��NmP	��aD�!P&����;W����K�MG�'�VO	FL(ɖ&�wW�U(�&�#��_���3ZN���PZ��k|T�;����[X�(�D�4��l���>%m��¸����`H��l�v�5>�rVP'sq�m�eDsy3bs_��밞W.Ov����D p�Oeá� �X(��Y��2�"��i(.�ˑ�4j{�#϶[aA�4�hr�&J��N��l�L��!'�׋��[��w�,�wb���\g�GO�����u�QM�Nې�z�h6r@�7��Z�ufc<��X� pg�>^g>�K"���`[�����	F>r����r����h������c��V��A8	i��8�Aߥ���mE�)�+�4U��M5@?~�n�G�:F���oj{��] F�Ds��"���9�{̞���L��|
��"�R
j��0���<�Y���0���PS*�
���V�`�E�K}���x��J_��@2�MNI�'|��U�R���?dH�-t|?\ �P(xi���?ݔZE{�N�}��YT�gQ�A5Dn�4o%�{�XJ��n�1�Ȏ��������� ����%<���h�m;�����J'����s�蟀��C�|ȃ�.;����׻���\��#��Й��r�����Ie՚wНM:���:Tvل�c;:�f�5�ryμ�9�O�~Ҋ��t ����w֠���
��٫(F��`��#.�n��C��o�frY^�f����m���L�����������+�'��<�/3[E*�O����8v9��F��a%S���u��L��+V	j�lV�u��ȣt}W�b�`�U]�8�F@z�A��d�l��f�54�i]��1��{�u�Q9���Y��hP�wa�����B���݁���{x��Є{d � �g��3�����v<6�#�6����xS`ҫ���Z�k�ϳ�"�o���Iyd���e��'�����D���L��0�y�L(�M��op�l�=C�,h�V����9�_'�Ie���64��&���	�݌�I��wTz���2,Y%�Ƀr��@�ޟ�h�����W�
�
������h���	�_}�"��$�Lggw��9�ܝ�Z�Mo�l#Z�-p�L	M�೼��(W�Ě��=��N�X�sy�5i��$�|D�4ҖKM���U��a-�8L`r>�wzw�n����1��ߑ�0p1��=a��*��a�C�1Lz���D��)xǼ�"Г/�$5u]����0M���Y��p�g!����e��, �� �����������EEYРB���D�g�i��W�5v�"��cw��7���uN[�"u3����s0�λ��#������A0�C�ı�pث}"Mc�?��@����	ɋ��t���>�{���{;o̷;��-���|� Z�gk�)s�����&�DJ}a��IVN���l�y�"�\UH����NM
�^sT�no\�������4��ݴC��t;�h��W6��J.@E<j��b9;zW�=m:Y�-R'�2��uW��ZI�����0"PLH
\D���A���u�\��M<�H���E Ih�h�ȱ��/��^�t檮�}��,�R�͔�>�����zmt�	D�&����"�����C�#���N:��o�э[c3N/�a,B���(���g/�62��m�p�ܭ��^��T��������?Ǟ~��~ <vH��SG���:HZ�ϝ�+H�;�0쬐��V��������\��><��hd6��mu�Ɩ@e��`YR@(q2�0����f#@�8���I"�ű����f�RT5wڔc�8zp���"�Ŀ2�
B�%�E+Z�T[��	����ӹ�%~��s}���y� �ȳ�%�I�E��7ua�J����d{nqe[^�Hʀ���<��!$�uw��*���F�`��J/Ni�B�X�����2�k���J�͍�0�<�gEfT�<�@��i�\���[��G?}FA�8=���7G�Q�*�C��t�P�k�^�8&հ Bc���ǡ��ƃƀ&������>΋�CR�w8���2���/h=T6b���,{:��?&���.���������0���N����R��<�)x�d��R�=$�K��0�J�ֈ���x�g���Nf�t���ä%@A<��� -s9F����-F+�"�7�.u�6���.�ω�f>�K�=콣� ���L��ɨ�L�L!3T��Y^�i��҆�}~���������`>�p�tB�0ϾsʜN�[����I�m�[,�Wc�����o�x���
���qys�|nJ6���#����-0�T���
w9��nٜ�Qs����9��F�]���7�ڝ�OtJU6�VI�Ψ�0��������ˀl��۪~�q�Vɶ��r�
o2�� ��G�����9l����D��*��A�)Ս�U����ėGQ�e5��ԥ���k��A�����N�d���ŰĎ�Y�_E�įYG=d&�u(G�?�O[�K�9-�oc}�q�̣�:��`�3q�R��C�j�j��v����a@4A���0��upV���>�.D���a�E�	 ��x�ͬ�����h�3��w�^�G����K�ʭ��A���An�eܝ,`:%w�K�aĶ*})ҥK�g���T ��hR����t�yͥStđ�_�~��m�o�:fDAd���)��XA*ߺB ���G��-wtʲe)�{a�!����1�#�����)_�'���Ɔ/���d���
w7�.�ֽ�_϶Fz���m]y$��,C;{�[t�4�>�������`�U��e�oD�?qR4�Tb�/� ���/x��Ԝ���gYfO�]z�e 8�K�)��QH�9��M5V��yR���Okަ^i���5����M�fռ"M���G4�.�(��+�X�3 �C�)�y�n�8���9�������KǞ�X�\l�y�>#4T W�C�����J���V���]�wvu K��������н��lHWf!c"�L�I���d�S��.C�$C 4��P�ہ�<�QC�^����qq4�M�k����nß-+��/f�?:�i���~�C�Jp���C�X�����x�ń�H�� e�L1SN�|�dK�]��w�3�4�m�HM&�#4��;q�Y�ع��a��u^���U��'�cYD����j���@*f���k�1U|e��x[�r�,5�S�a�%���q��!�B��/teE.-��g%� ����ş���=��<��etu�7l(��nH��fR>]n�ƅ�Qc�|����x_c�l��:�4��~���s�p�2��b�Mj	�^���8^���,#*���QK��~ת����
#��Fh���Z�$N�M-;�:��Ǆ�"��{���,L�{^��&6 #�C��C������Wb젟R���>�:{�d�x�R��8���U�X�uZOnĔEXb3ZCb�367�518j��\�``a�1
���u��t�=;E�RR5ؽ�-P�/;9|���9�(�4�����l��~���p�	�>�T�ھ_�+'����I��W!y�G4�� ����� �������6M��P���QFJ%-�ӱ��U���ei�Y>����.��u��e��id:(��
vo��ǕGJ�{�������gO�{)������W4ĘZ����!���5�h�}"���^�Kذ������e)����e�3`w8`��!��>���U�Dw� 3��JqD�>[��J^8j=Y%�B.ל���9�>���:��q����-~�/3@��=��%CI�"�H��૑[�j��f�&�ľH�b L���bhm��e6v������Bꅺ��^�
�Q��������"pU��z������$<����0�'���P[J��8�Dv�e��(޴9OJq;Xk�gc�̴�������OB4�̳4�6צ/f��D�0���H�U��EЁ7@|e�B��Ȏ8�>)�i��B�v�����G��;}Z$p�������kA���k
 �Y����U�g���ng��n"����~�}��2�9�G2�g��1�J>�;lEWq)�<a�&��F����3�u��t�^��c$&b�лzS�U����K�ԦDE�N��Z7�ÇlX�gA�J}�x}4���^>�����ȮZ��uK3xΙ���T.�K��G4�a;$��$�* ���ǰ;zE����]UHL��-�?�=l8��o��q�ը�ۅ���U@���X��b���d�ɹ�C���?�/�Wd��؋����)�j�n�7H��P�u�;6@���>R�W�O���ͳ��AK>>d�u�:!�`�M4�+�w� [u�P�la�������?��sqw��
4ETK�,A�~���W�A�c"/�Ї��.NRq��z�hu��uX��$�00�	��,g^1����� 6�B*�N�G+��.�w!#�3Zp,�8q�0+؁O�s���p��jPk�&y�ja�{����P�F��Fw�D��`�	��SH�U����<���_��3(IP|ڡcI?@W�ǃȪ�-�*��p�7ĸ��+o
�Tf���.� �'l� ![���]�L����_]2����F����Y�lg��H1��)N��3�/T�ؖ}����@b��Y3O�G>���'�t*3?�X�h�H��]}�-T�zq�xiT��az��`l�p-r��-߭�"��	Wbí�?�ü��!Z�R����s��:�8ޙ�N�t���3Ң[�f#�<�@n����	�7|1��-H�P߭�^%��y���ݿ ��5�c��7nU
T@�7%.�=�$#�۪o>�Crp���o�dR��
ª�4��LS����:��K��	�=h��QFP��� �B �jG�Ԫ�H�gOJ-��F0''uTK���A�w��`��?�2�kŇJtbfY΅es��)^z�4,'�轏�T'�=.8�����>�/�.��}�a��b0(H�8;磈Ma�9��[�T
�����;>z��,
�좜�vW�c��	�K0)�G�1]F���xA_k�:e1��F�+��F� ����*���sbQ�d��M�Zs�Z��A�����Z������r>p�ɹ��)$�>0������[���6ƭ$��.$@"��2l+Ʀ
�ۂאҙ�(�p$v�|�؁���
�{�tY���\$g��x����G%=Z�p��S��͒�9M��d�M�YԂ�jF�0��I���RD���M>.�[	ٚ�E
���i�ﭱH�`j`��>u�Э�.q1��E�65p�{��/{���@N��1Z%iN��I�l���u�>e��!�j�>O+(:e�:OĮ�li;�bMM�g�B�ݜ��ZQ��Ͳ���>C�it�t�}~6���{Q*I�xg`5�;�H�~���k�7%�v�ꉼ�>*ߚb�-�z(�mL�T�1�o*� 9*�5:��7��|�S9^�2�"�E��:{���¨pI�s�Ϳ��8�s����e��}����<�Q�0z�-/6��"U6��h��!�u���<��\:�~���d_Q�����6�����ÛG4y�*��q�_T��{���Bt�`��.�~��Mw�d���[��u|� �e&��,�����w�9� {�{�&|@�A,�]�b��'��8S��f�h�_�P�~�XI^[�/j�oc�s�=Q2�b��f{�
#Hj�w�^]J����G��`�o��M���O�t������^V��"u!��$���L����W�~�聶'}"3�PI����\�%�Λ�!��:6�{v�z#�߈�	L�}+��t�MZ����*
�3�"���ʅ������A�����
z����%���5�|O�LK�4��	m?j��ی �S5ૼtx�ԟjQ"�q:�q6]*g벴J�S�U={^Z@�P'έ%�ns��D�>I��Np9I�K�	�<x�йj�����i����#v���=o��~&AcLT�±�E�f:��}<Y�@΋NDs����s�zO���$�-z,m:�w͠�q�P-�L}'>>�[�j�Zt���A�<�������f �)��¬ڻ����Q'�����@sY>>G�3�]��ע�e����7��~� w�Pa�U7��ջU��Lj~ۚ^�����~{��m+�[`��;�]EaOcʏ����{d� 6\ڗ����q��z��̥�6R!��C�Ύ6�*�&�j��<w���w�#X��5j�B�q9���|n�Z��nKE��BU%�GE�C���!��Ƅ2�ŇN�ǂ�TP��^V����ޮ�tJC�:2�M�Ů�qq�a;e� e��y�9�V�Ƃ5I���d�t��~kU�ѷ�5�W�KG��ў�_����_᰻���mD�M�X�$tuǭ��3��nĲ
���qSd���j�%�=�6���ut�b�X��8GD�0��%o�Fn���N����G� ��[2XPR�N2�XC=D��E����ŕ9Խ]u�L��!���А��7����r������_�I�$���Imf@��_i��	�oiA#��od��K�J��=�v�s����ϻ�)��P )q`��x4��M�k:������)/�~AёF���!O�luI]&u�Kh�D< U.,�X$�j��H��X-����o��>>���
GR�5����*�?�c.�(R�N.��"?Y���Z5�^,%Q�Mh
�4�s��_�����/��S�ӀFJ
��z��z�C���0r�U
�
PE�Z�z��ؚc������X`���a�ǂ8�IY���LTL~=��K�̓���ސu] �to��/���uN��-�`���aD�dR�2����=���LS��p�n���l����-���M���'�bu�n��^Ȯ����
��]:�F�M�]�C��R�p>G�p���*y7?��T~����X��r��9�Y�n~��P.�U'� ��/oF�_(�)5+H�㣂~
^~r�x��:R»����9�7ctC����I8�}BPP�ec8������p�|8B�x�f8��zi"�_{YŢNS~[�QD�R�)$�y���X���\٢�ׇ�~1s��&��0oSX�0�\�[�>������K���Ӹ���J�ؿڵ\�R#�*o[��n�_:ǁ������=��	>ٝ��S�?.�cSS�4K���b�#g��>$�O@6Ei���0yF�,�v���0uJ_]��
0��ą�[�x�=�WB��������e�D7_����(o��X_[�}[_7Lx�7�ha?�ab�����II=���r�rޝU�y<A����-b��;՛h?Q��
�"Sݱ��Z���0O`zA�~�0~�3��$d�!����J7mZ���V��ϰ��,�Y�{������Ý����l�ƭ�o�_��z^�3��ۀT��}�ߌ�T qؑ��A+�[���+O�%?�e�{����׿�&���.�a���	�g�Q����{��1Ĉ%S�U�8��=@cw�ߑ�oOw�*,hW�]�	�|�6� �Y�����F��x��%��A�{�c�f���0W��'�HCQ�s"��vX�º�5�و�3��D|a��M����L��8�j>J����[ͯS,�'#QAfa���%	"|�U?�.�d��Ɋ|�Y�P�݇#��bQ/��mSv@�*���+� K�wE
�Q>C�v��k��.\be�&�t�Sj�dK�����N�6sj���c���3T��޽[��>��>���.%%��:�_�䁚��_����&<'��[�У�j���3	���4��@�mm���]�ۈi�������p[�}��J!�#�ą+e#e���J���L�k�HL�1��W����7�K
nb\���4'DZ�4ew`\D$���u�R�s�Yc�0Ϛ#?�}��e�gJ6��
���0p�ӌR�� �ST0��wl96vK��~�b�hy�"�y	����	xqa'D�Dn�W���!��J����=N�Phj�<�:$��nJ4
F��*m:z�JLu��~"�vS���8�b*��t��J�`�V6*���Xf����<Rn����v"��<�4=�����j�\������z:�]����#�^�����7C'���P�/X,% �5rd�����oLtP{���o��IN|%?,�ӌ㬻�97-���c�f���o�@@T[��;�����)xjI5��0��D*{Q�P��0���O[�ٰ���������/B�ꤐ��jJ>��.Nj��m?1m�_�v��^B/��+� &h yC��P�R�$�Z�E��t��
Q���:��c+�0a
W����7�y�F�ysb.�ͨ"8��a��R�]fF�ígʬ�}�\�\�m��c�t�)J���y)j�����4'$k'Q��o��� &+��R�������Y���r�Qx%ն���{�C_af3��L�}�3q��RIv� ���^PR�����M���j3�
�aK+�ށA\�_w�j���op��nwB��yϊ	n���x�D��^�G�U���-��_�i:�cX!�^�Q��Ӈ��`! 3�S8�G���I��,>�e�'j�cFr���zZU?�P�D���z��)�Ǻ��'&C8��]+��\ �+,���\ҡ`�PI�oW�p��$s �Zz2L�E�Ł�M��,J�yd�o����5��*�=nT�f�V@N/�p\��H�h܄W���8�p�h��)����� L�̝bI`hVYg�l���)Тd�7�-��6�$��,e	��yl�~�F&Sv���f�	+���#z�5���S#x�����Fu:�ߚ����`,�T*\�k���}���<�m�u%�������Ҝ�Jg��*�K?:~�.w{���;�<��on�uui���ޢ�z�Ugs�&�YÕ�@n��M�g�	(�V���c�	�-��M�὞�<���,gG�)�(j��˔Hp��	�D���H]9�>�7�����B7��"�M�*p�Z��[Br�O�/S4GT0�03;I�O�+qo�����;��%R�ړ;���lV��p�5'XҜw�k���$��ň�+1&KS��|"X�A*���Z��[Ɉ(z�n��&�/�b�roO+�}os�Xv ��+4����k������Y6X{�Z���^`M*����&���4�Oſ�F����	L�O0�mF!D�F�_n�[��h n�$�n6g�FH&R.�ã���4��ߘ�q�JLW�5в#*������r�Ţ.wV�u ��:�;�錼�-W��H�}���_�t��<Ie�qIX`6X�apR���RqA�-&��*�bg19��c[�a��f��A�O�C/"M��5��m_{w�wtE��E@h���Z����M�3��-eEK�b4�K7����?�s-;��8�	���}�R�_�� v�n�#9���M�HtƟ{��7dq��D-��C�~�q���Ź_����*rČc��?�<�����C/�D�:Y]����ME���G�0c������Q�����J��P�&�:�Fܨ� �6���Bk�z5�J8�g!�%����;H�H�n8���(�^[�66��}|͑�Ug~p����lOfJ�ppT醴~��s�>,z�1�@�=�
��(NB����
��p���j�	"��\��sn����1��Mi���h�����=[%Mn�|T����zT)xD4�=��(I5L�� ک��Np{+���f�4��$�#c  ��l��SԴ�E@q�xw|L4�hS�PƋ[@���Z1� e������-��?%����FJq�/,���O,"��-��K� �҅���.�Og�0y��[����_�K+݀�N�sT��z<sƆ� ���ܵ�^| *4p��V��6We_�k��
e�hIl&�0�N]��	�q}u\���bq
D���ɌU ѹ�7Ye�lh�t�W�6*�O�Dr��ދ��ʔ�����	d�����p^��/m��9%��ު)����Z=T��G�G�1�u^�#����)�<ٖ�ǟ�!Zrt>��9��i��+��i[h���z�����2��Z��	w\�Y��4s����M}���5�x�|Њ��LnC4�ܩ7��΃�+G���KA����ŧf�Z������(��u���<��k��1��o}?��Ɂ�؍)m�~�9p�є�=԰+(��qÊx�������)���XϜe���!>�Q�������:�M�1��Y  ���g��Yǐ�6U��ए�'C�İW�$���ws���J���[����eu�M�p�0Lc����l,��M6Y͐r�ϳ�Z�ů����FfC�l�{��U��j
�\�1y(���oN"������,n�;%m��4�[zp��/����W�Q��U�s���` E#�B1���A=����=�#���H�#���2�Z���m$����]�����n��UWz@�{�оP����?�����T��>
��Ep��D4S^2O�(*��z@��uڢ���O��|�sT�UZ4{�&�r ��� �w�ώu�e <_In���"0n⾿�x�4�+�	َ9�Ν��ɗ�#���R��ҒR:�<����Sh�>��g�^krR����.f���c��(ɻ��"�ы�:"��B8�zЩ�3ң�<4'��A���V?R���/�t���X\�x/�]W>)̭�i��(/N�e���;-^�:.r���i1)���<���g��JM2^����X
�[h!ȡ��س�<�
~-~.�Σ<�]L�_�mb����,�~���K�)-Æo�˚�@|���-]���Q��Yd�pZU�(�ⷷL�&v���TX�X�C��L��Sۊ�5��7��O��!WT��H\3w�_G=�ؙ���5Hzrc��<�?����rj8x`)z�����}|�NK����{2�^��pKa!f�c���oc.G(�)�Jz���Z��W+ݖ�z���*��a֚�����X�:����b+8|�]Xv4�:0���lּ-(���<-��e�F��0�+��AF0T�=�Rp"��	]������CG/�7,����w[�!��%7���mJ��t�p$��a؉���,b����`3y(����d����v%�!�w�O��w�O����^t�uY�nwS��x�/&x���~f��J�~���6� ��&x�1L���	&{���
^AJR��Y��< � Mz�]j��ѱ$�-�	�hs-S�V��e'�<&n"~Z�?��1u"KhoMU�("3!��i���ڠ�^�C��Yw��	�R�#=4���U4u�Wlp/�k�����u���x�"��U�����l�t��D�5�
�i�~]5O�kY���33gK��;�,��s6�]��F h��s�A���K�g^���V�h"�?n�6՜jE3٥�k�n��Y����}g�4��pYy�{	��luB�?�ё�9���WHy+�ż͢�N�}HtS/�~~(<<� 2&��Id�%��� Qa�i�v܎�8�j��XY�Q��9���%���������c[	j^�.�a\��S��D`�+܃�J�;�q��p������7��;w�"��%$t[�2��Pg\?Ԇ��¤�$Q4���v�L1xUD��MY�/�"'����0��o�����S�N���Ȩr]�7��c'��#�� ��3-����WT9��MJC���R���Q��q�9y*%:g�C��G�s��#)q"�p.�_�~���;	E��* �,�j#�6TT������>N'�8b��{��<%�[��fZ�q�4�z�.I����4�$gwf3pT�L2����6.��6��~ZQ"4�.�I퍚C�pd����Eh��g�����P���:�	�CY�d��M�{4�A��Ï��c�Mlvc =�������E�^����k�[-$VS��hn��e�0���X#��|D�q��q �έ_�f .�q�s,]��h�n�
nC�C��s��=�30�q>`�H1�� �0*L�G.՝�f��:.�L��Ŗ
��Px�]����,pk���y�l8�Il�ym�1�1̬;FMj$�1����2��%/�˨)����R��w��D=+u��6��{�mX��Z>�@�����ve�r��Ñ͠ Hű3�k�IZ�T36D�0�������Ŋ�nQo�������`��YBn@��C\�62fR7�~B�:�&`���洐�h`�������A�n���_������94y��L#J}�g?>E󀀯��x������f�f��l{iK�7uS�*S5��]��]>+(T�ᩔU��	u�\�&���y�; H�)2��S?��l�w*�JݜC7C}����E�����Z��c"Dv榍�>g�g�"9��� ?>p�b���tN�f�����í�~�]� ����Z�����~��]�_-/��f��z��gpb��3�j�t!aڀ=.���c';��������#~u%e�■���$��V��=����^S�/Y�x>7^g�/������R+�w�b���'[�5��V��5$�޹�X�]v��7Lx�+N n��cQaǒ|b���1�E��D�}��N���$�m�ti �o�8��<�@��6�+�wr (]��c"il���b������-ol�s�	�8�J(` % ���[W�|Ԇ"�C��0yճ��;!�`uqh�/rr�0�o{}g���z/�]�S�7�������an2h:��:E\x�4��Y��O=f������.
�Y���r��=�Z�����d��%��e��݉@�5���D"MC�[D� �M9��VhW��ب(H����sL��n�#e^dn���U^]�8/��V��Y�6�˂\'S@���8!a�,dsd���N(�K��pE�胱-HVC���/��):�<�(�E_je�,�����D�!�@�F���Q�Q�V\���A)�asP;���}�D��.l�^�S!�{�����?���8m�D�;��0�qb-�F��k�l��X��͋~��۠�3f����i=�u�)G�Y4H%�����(�[j��> V+у筼���[�5�)j����p�tߛm�I4�mGP@�w;��ۗЭѰCNVc"Ġ�����uM�O#Gt�s�'6��a��]}�,��lO����?.��7�����giv�@�NyX���D�v�";�^~��ܺ���!v�~���������l����@/J�.�kЊ��كH�UI^��lX'�%����a{Iu�R�m�7����&:�v��R�3Y��@5�R`p�>|�g5i�N^�!*�B����'�h��Sv�o�����7��p����a��b�?��#�,d��4[=��'h�`Ǹ!c'���_5dկ?澂�i�����r�lі��
���\?��0Mk��$w,6��Y�Ӭc�8}~Un����V����z:�x��u�#t ]�6o���]���"ę�<>;��/ �S�h�Ȥ�u�%3W@�;:���D�RhR�'B�^cwf�/�f�f�S���3>Ā��2I+N�0�� 
����N�]0n������3$����|Py\)��b-�91JkLN��q�
^*p���|��9k�y8������E�R�[<G�q��f.�Pw]��D۱�Y���ʣ��	 .��u~�W���`|�`�#�:{�gP���Q����,�]�*�(������޾�߭�> ��Q��/l�BЩ�ۏ���ls%zlh	��J0�*_;c��F�P�<[ß&cI2�K՗l�����r�a�;�����}(�A^�� hN���y)�ϩ��������3��ӂyNZa��`D�X ��M��t�)�A��%�ь��6���Ջ�B��"��(�A�7�df�����$i�Q� �����v�ċ��B  ��S�|�i������xKS?V`|�:�����;�,	�qW������,Qe�*v�ng���N�F�0����SBd;ૉ>��F�tg��Cm���2)j��4N���[e&z�Zڽ����=­��c}ŝG�)��a=ݕ+�0����ԄYy]���ݔ�hR�1�`0���6N���bwp�2(�����W�h�=}�f!s�j
\���Nhk� ⏆��!�Q��?c�l
C
,FW� 4m'�H��z��s$L���ݛ�T�hz��K�����a?��IHъ�*$�E������şU�_;��X	��	>�6��{�bh�T_��W�����刹�פ?���i0�H�Մ�mbL����iY�ڽ<jX�r��D<�7���1��H�՚�Է����y��b
���6$�"R��ބh��tg��k�������:�#�q�g�a2�e��Yx�����|�0.�nҵVΉʍ�gՄ)2O叚�J�UH�) th��LJ�x/��-�sv����� ��Fҭ���:5�!e�545��%{%H실"���z\Y5�"��$5��U��ڸ3�o���>���n�k3�=TM`t"5��Y烮I��ut��E��x�'����CI�@$�T���'c]�t)N'''�<���Y�o9��M��}��������*'�I�%�&�Rb�/��7����}mO�{��RJnh/���ۅvc�<�J!Un#d+Y�^�G��.-�Pe���Z���:D߀?�!A� ������qǻ�&��rp��0�'�$K:�KiC����1����rVs�[Nm�u���n$r��#)�����N��e�T��>W��Vb&�5� �p좂S �Z�둜.;�m�k!���o����Ltpd�)�e8��9]7���j%'VZ��/�&��}#c������\�תͮcΆ?{�a�jPr��˛���T� Ro�1��O"5.%ܙI�?���oo���h�z^`h����IE7�g/d]��x9��?�
����F�B❘���%�T_�{���bX���汦���k��(=�6�۠p_�ޮ�Bot���)z3�_
�#��N
,�PC��	�Ze'�5C��m	�c�u��+�u���VyW*=x�����i���9N7�e�d�}�yL�]��?򁮰N��n$���9�k}���?�;��B)C��Oѳ
����
�
�X��3��2ҼлY��u1����j[�d��̠�����/�ֈ�GHNohi���?S����龊^]�)����S�ގ]��7b�	���!�ڣ�A��b9���gjjq���.��1{�?�V�9�x�Sw�H2.�V[���㏂<�i���P'>&����]��#�Nl5m�=kf�r�+g�Qq�܃;le��O��jg�r~�v�� �MNOG�@�Ö�P���/-��/�Z��nh�� W�b*���i_R!��B�S�P	��U~l`TA�TE�� qk��I��hT�	��I�p[�I��V����Ú�ܕv��@���ʱ1p<������k|�Z�TY�9l|�J#'�8r�l1���,�Sn�?]�]:%���Fc8��ل�D�ŧ^���:��'W5����K"������pw��53�訅e o�-֐¦tЍQ���w��v E^ʻ��� ����������
��h�I�ށ&�X����.X�f�֛O�)��9����^�)\���/�"}-�J����)�DB?:�{�sm��8��N���E��Ec�iQ=�z�����5ϋ�N�Vß�y����(������ѕuz��P�;�¬I|�tu˂.�C�]+E����(>��-
�{��hm��f�;O�cg����>��_�D� .YFJ?���4B���4q���$DB�Qz��T��|�A����Y��$��&�1���}��R��$U�L���xya��IKf,%��x�0[�|�zHE��mE\������=d�r@C2r�'�t��B�弔y�Z%��+�x4'U�zs)g8T��Ɇ8��������d1#3cyu�b7*b�m*�E8���zp�5�p�Lq��/����(��B�t1�-�ȵٙ~�v-h�8��?X��L�V���sC��sQ�m4��a�$4�z�󪺽7]�)ǀ:d�#�pK�(�@t߶\Pxz,&��H�m�}7c\��=;��w���L�d��,zl��TՃ��E�e+`3*�`6�ČL�k��Y����6�N˹�6����\��٥7��1a<�L���?	��A��[�������qO#TA{V3� ��%�$�/_���άN���HRJu��ҷ��w���a���%(�Thop�:gx���Cg�k�bÛ��b��"�"n۲�*�<i.��ϧ"�s]Ϙ���sr���i|Z��V�H�S� �]���ƺ<� `�P�O�R�>-�7�J��N�C����1%���Ky�L���\�t�X�D�Z=7����K+ѹ�A��s.6��`��o�;�E�=���� ���?��C�@�X��� N"�����\44S}��0� f��w��cj_u8h��@<�;�?�D�6%>?:��/ʦA�?�Rs��ݮ_���&p�;�L�,O'�=�ש�k���iʏ���DD��Ѕ���*�� 2HB�ST#E���J����g���x`�Z�V��̼� �f\�[�#D�=�4�u5��� :.��l�UL�ʑ�s�C�����׿�As�^�P1���>�D��!�J����7�H����~׸�z2e�#�V@�#&�	N�@bʝx�Yۂ8`�*c9��jVmI�e����(,���� �4� ��n�,iZ�'�m2���(��zjd�H�F�hj'jWU`)ŵ�L��sl<�[p!?�\>K�Z� ���^i��A���������l���R��ݙc�����2�����5���u��Z�"@�f9@��=����G������[��^��$O;�ѧ�l`��F`E�����Ca�9���6��vi���O[�9�}�q��m�sc��So�D��ShV@�3h1u{�zW�޸�Z��-&� ��k�r��32"�	����D)��=T6�-A�&?8�WgE���c,F������#��Z����H�ȁ���qy��BKܝ�u�Yɏ5�]�����t�̋�Y;ƫ5|՟�n�Kǻ��D�G�
�>w�Ϭ��^g(`��0��=�j��
��WL�dr&?���.E�ա蟆ս�{+�W��E3w<�	W/�O�^��9Eo�E0�&� Ѭh����cl�MȮ!����Ů[�	��Uz�ο������д�O�,���w�TJ����f@=ey�h�[v�$:m2*�k�kQ�@� �*[�z��^>�C�W�e��Y 뻘?�M덣�±+T���9L�iX���%3���GS��&��`.�y-μW\@�tq�E�I=��K���8w\{�/�5�B��#�t1(#v�'�F}���F������� �?E�
�n�1��*>��"P�G�ŅfT]��!��b�Y6?�u˞�m��>	��	�����I�<md3չu�(�~G��Q��Cvr�����8�ԙ�<[a�w5�/h��K�~I�~��fpm�^WgG���8�|#^�U8�����tb6
���W��	�s�PG��FCFF��^514,U�Ą�Xo�g���)�ɢ���:(�N��q���*/��*ͻ�g�k-m)�����w�N�m��e{��U��m���_��h^�ḵ�}�@���k�L���`�1M���vK���G<�����"�'�Υ��@�[b��sc���m�H1�3eQ��N7.�|��"�Y`0#�{P��و�M?OQ����!B	0��2V/ 0C��Z�v���:�ы}�褃|��5N�I���\����*��C~_�A����n*Ӵ���Z����XbD�,c�n���x?�#��ހ�必��|^�{��� R�\��|������@H+��WĤ�C`�}����܇��c�}�u�-7)޴��]9ӆ��C�M��3��w���z��5�n׽�w�)l9F?�%�:7�ڶq�Ytޛ�,c#�+��v������-�)ֲ�L?���:��wA��������r�\����%��p�EH6
g�"f��6�b�ԅ�_�����x�
���*!ͼš�;ߣRt���C��#��8�T�V<9�(G8քi��F��<�P[�!&�I輧n����O��{{?%�f�Q=A�ٮM��
'�-���_�f�@�(C*�9��Pi����fY� ��~�9���V��iLq_�3�ÇA����̻�'=�	�`Ҟ���9�;A'����Ҏ9�H{*&���-O�Q��ٖ����G0���]����2f��s�j�;5�z�B�0�pXw��Է
�f`��!J[/J���:*���hI�3�\��%J��2����o�H<��(dPVbM7���������4�*hu���!�@�?�3;Y1��Z�(��� �3`�GMX5fYK͐���6�qN�z�w�D��z2�(]ׄ��W�;�� F�����V~M#��~����ι���71:�P��ܤAY��ǅ����4�<�_������Gq�Ct�c�{���ƛ��r����H���)�vc,v�{ F��Y`��'��q�ۊW��"��������ݬ���0�����OE�v�;�~Z/y
[<g0�'B1J��?��������6i�vZ`�?��U|RC� Z�o<%�x�Z!G���R���9�s5�geA��f�bʎ�//JyV�W����f��U��_� ��H���K$��-iÁJ"�Q��X��| �w��#yHYZc�����cm^�ٵ���~�>+0i��2V�Va�G欞�WUmJB ׹2g�nȘ�En�!��h*�v04/�r�]C�[�t��rz�H_|��fi�]x;��7�z�$�C��.u�R>��o	Ѹ�y��v�qW,@�H{��������I#�D����o|�+^{�&k�Ӿ���>�8�ο�x�ʗm�� ���>���?u�z���e�8VH�͋�r���:�:x���n�>�!���a9�V�a�����/��޳{S ������|յrJQ��NR��:��ڥ06W4a���� *��ƴS����L�X�]p����,f7,�ǔ���O�R�f&�(���h�(q��*�gH��aC|��'%������wU��Ot@D]��*���y�w�""~������揆3Ar���1`���m@zh�T��-�	v�3�2t���ì- ��u�ݷ.�=Vl��ԋװ�|u}_Zq҂!����#�E g-Ӵ��K�R�]��X!8�L��T=�޻�C�'��0l:�TN�ﾨ�i���y]���纲�[�v�������;��{0k���;ŭm2����\�բ����&�X�����JD�ɨ���\%-��lX����0+�}	Y{��#M��S-�8�]G��s�gB��C��`5���`{�H�v8U�b��{�y�U���&��1[��������EN��x�&&N`r?l$
7��S�P�� 2
���kף�-%�4#Q��Mf`�
1�C
+�C�$��^��(O���w�����z#r<v���ކ`y����|zUՉ<�g�}��R��eS�pv٘	�P!Z�YR�	��ն	�:/�&t��<-c�;�NZ�3v��
�����UR
�AGd�ak.�&=�&�+�&!!{��X�Ur������Re��Χp�G7G��>흧����nh�/i�g��1nN�/C��Pd����w�Z��(����w�t򏾭PX����Tf*�xMtyR���@�*\���Jǒ�>�g���Z�᮪�lє���d���(̸(AЀ��7
5ϥ��cI���Jޗ~F!9�w�P-+@�f-�SW�.п�YD�N%��f�ru����i��M�B��WWN}�$�׬d��9�]H�<�g�K�z���l�RgE=�6놾[�)?iH*Iv'�⤼<�@�	p�~�%���1���'8E�Q���C�{ʮ�K�����ؖ�kJ#_'< MV��wVb�J��a�go��ė����(��&�f��{zy>�~�,2ź���d)�޼n)�'lJ�\�#�oc�)X���E�sK�Z�|s�I��_<»�7r��}BW�u�!�#�;ΞR�鲯��n�����5Q��
�I�	2�ɉ#G���(����WD��F�(��s�9�4Ͽ�t��9n������n�/���^�&qBl�3J�R5Au�ȣ2 ���9�"���uU�C��pw�5M�ԩ�DK�u�(�</4`�M	̠�����ڱE��-��?8h=�6fT�@"8�cƮ�4{�>�d�%�")z�q�pK�2RF�6Y�mX�в��+}�J�r��F���+]��35�1�SH�JFx��L0�)��1�PY��G��ف6�[q��_�D����R�%Ȉf�$�<�?@8_u�Ŗ���f¼:��4�}��_��SwWzɌ����ADFqHR����
�����8lzc�	��V&������[B z89.�H��c��W!�(m�r���>�;/K���aE0�.r�}�����"�Dx� �
?a����R34A��|�/n$k{�j(�Ēˈ "_almϰ;;�B^UHƀ�~&r�R}V�Q|X���e��_w��&�V�ʜT8�� 7� �G��\��U�E��v�S)H�'6�5+
���q�ۍ{l�!B�"E&���Cf9�e�[c����B���[�҄|Tn���N!Y
v·ƩN��� ��:�h3�~(]�J=�� ��N�=bd���)=���#�38a1za*�a�i�B��97�L\�S�S/�|w�.n�����Z��9�n^O��J �_�%�~&IW��~T|�@(�$�+�<�G��t;;T���+瘦W��s��(�[u@{���w��U]�&2r}�<���Ꭽʚ�Z)b��6��� ������YNr��D�d�dl�X���x��cZ������͵o��<ft�#=��V� 1���0��O���
ˍL�]bI�K��i(�@2Wq��e���I�L���[%�+�;����ig��*ɜ�13�be�?�k
�>�g!��;��nw8O7�)m���p%&�CLs*���^	xL,Ѐ� 3ù�[M}��7P��Mv���$�8�E�M�A��_,~���4�e��QB)s�^f��'AV�o³��r�̞>��h�'���t�O���`a@�!ë�"k�V�6q1̣L;j�rK������@0]p��:ݓ�A~���k�e��O�$.��䁓c�E%��:����\�_g{r�WW#� h�S*:=8��F�t��9�+Ѱ�()�4��)E�~lp��;1�(z��XuA!v�[�"��5dp��2�Q�hŔ���0�����K�nd��+�����1�}����N�l��x��KU���F4�P{�������
"�v��~��h���֯�̶�$P�Վ���k���Ħd��֪���gg��,�yנt��$)������O�V�/��G�PΆ!��:J��?R�w:~G�(�Q�{�ClVbE���'�y�"��� ��yC�!L���b/�m�
�5&��'���VCؕ��L68ax�yY��ܛ�؛=�"�ؖ�c,HU��*�:_�����oD)YZ�5 ]�] ^o�$�.sC��i܎=pӾs�����Q |���>,�«�]8({�b�!G���%u0� ��h)�ZV|�y�o��� ��闘8�\X�<���i/S�g�|5Dϙ��ײfa��:</�-E��}wH�ϭ��E����Y%��v��E2����d�����pG��H�w	1�ݷ|4:�ѭ�8ӓ�45�����w����������J~�+�bQHH\=�D���ʷD�h���Z�1�u�"Y_Z�w��>�s��������Nm�,R���yr2���WIR��6ϟ}f����>B�n��x[k'Nr�i}<���/A�2���Z=��\��0��K�W�"όRQOEa��y۷/���ˠW� 8G����!��cR7{rV/�N�I��?�;to1���K_=����_�4���ݽ!�/�P��י���4#Y2�|� �s�y���p��N�ؙ�dB�;l�`��rl�@�X]�&8ԡT׺Z�;�H�>¼id��x$"��T�1)�����?��}��`�p-���ѷr��t��cfg�I,[���{���<�"�����J̇��W��c�����/i��Y˪��#I.��Զ�4ˣ�?�z
�!*���ka��t(KTE�C 	�?Bv�
S|b�"��?�PXH��蘟���to�g�'��B�HC4ٍ���)�7�	5�v�d?U�bw-4!��1.�r遈l{K߼�}iK"(��ݡ��*�'-�C�{�_�<Q�>��Ys5!�{3�dm�#����%�8�I>7<K�Y�϶��M����
-蓶���)�A{Z<���Of��ț����".�5����̦���.23�E��oy΀q�ϟ�6L®������cc�:u����p��$�,�7<j�O��Ȅ��em��Hr�e�5[�I��^�*�e�����Ҍr�S����2���>&uzs�n@��w��մ�lZ]�a���4\(h��}k�'M%<��O��iu���)�'�엝�_jK��5Pi���z�7�gF_��T��ˉk_4�g��~̥0��[+�)@�?]���7Y�Ñ�I>^�r�s>�3�j��(�_�{�Vo%c����0 JG��5�,�
`Pmpy ���g����M3'7x-݆-��)koAT	'��ɳ�zT��#{�'m�(V)��:+?o豟/��Hr���a��PGςE֩e!��eir���R����V�=#���h��$湛^V�v��Yj�Ķ��G�5M8ʰ)!�IH�`�@� ��aMV-;�$T��i�xy�;c���a7����n��+��R*��M���l=�� z51����GT��J_x`s��A2'ވ��I�
�6�]TPv�	���cp�bBټ�[�+���񜊄�}�e�H�eLX��a��Z�k����O�+��^���5G�y��]�r�g��Q�:�t���Hg4���Ro��Wh����W�~b�}��}�*MD+{A(x�Or��b�3QH�P�_|!�	�>G���O�Y4
�1�GT��c�#d�c����%֋��;z�I�g�
�%��x����c��F{�q��/n����G���l��ðm��f�
	@Ge3�ì�c)B��aTXv��-?X���-����1'B���F���/���Kx�����gL�)�
rO��1�h�l!����a�n�/Z-��G3�������[�0��p�ʪ˯(d��56uJ+K�'���4+�ȸ1�:���⨮z��!���/n>�^ �J:�G��Ji��F�eʒX��"�yZwyy�^��fĐzR�Kh�X�ss�:"Z؎���R�w�A�_��AtK�1�5��ɹ�#Q�r
#�z.���Εq��`�p����!�'r����v��� f���%0��_?zC���@�9� �]3����.Hgħ����@PO4{	z��N5���B� �.�6�'>Gm���hZl��7853��%y��`ϓ�Ú�k�5k����;��j�2yN'HSP��� ��A��H���_T&��t�/�\>�����r���H�I��L�n`Ѩ��n:��w ��Y����SжY�w|�s��!��}���	�����Ro�|قZySO����
���3 ��O�^r�23i�TUC*����:"UH���bZ���	b�?g�%Vk<�*��c�����mL��'*u�	4 �"K�gGt�)��꣒��7��Z�z�M�U|�V{�t
:�]c�N K������9_b�PE�Ik�I~r�;L.Zh��LE�\i|��4�q�D��:�UB?�"�%��!AG��$'�������oG��"D�m"63+m��%�������w鮌�q닽[y�m�G"�,!�(ڄt��6��m$�@?&�:�0�lS�.Z�+͞8���Vi=�#�@��҇}EI���C��Y�W�EF�P�Ź�a{ů�l����dW��)W�d�������wwPӼ50���I
�^`%5�5#C�7��2眩t_(�Y�m�!=gB���8@������ 5҈��"��Y6p��Q@	��2㴐eI�8`�1�7V��1����b�:ye�+���7 �_��6Pѳ�F�Y#��!/zCj�����ZiB~��wp�y��v4 1k��ʀ��՞E�1�2^ܻ������e5���ōu��%����ܟ�>�	��Ǵ�v���C��X��m�b�-2�0{TQ�_>�w(�jw�ܾ�2妹<���|�K&�!1���}I�����{�3��,X%�>��^�E6D[��Ȍ����/�G��^w�R:����)�Y��O���v0�3N���';����.ڕK.��\�kҨ�5������io�C Б�GNM�|�����%��u�o~�a�w���`Pp���W>�g蝒Q�AO%�)	��7�t,e���9T4�ib�*|p��YѸ�8]�mz^[�<*`,��M�䊢��%gU����#�MM^��6���b!�N�I�ϒF�s�m��u�K�yP��6/CŰ5�`�ߊ9����n���n��_��f+ҝ噯H����/��%Kޜv%|�A��*�`���y���s>�Ml�t�?D_������^5���7.?����7�I�=k��▽����"{����m�.:
i�*��iy{�Y�o�����Kc�qR"���&��v,�!	Do<Eޯ��"^����Q��5- )�_c;�-	i�dv竑}���d5NNP'^����y]	B�P4�`�cQl,��8�}�����������ڤF��%j��T� �3���Yh�W�~ٞ^���`?�������P�ZX�7������e�uRZ�@��x@�����?g��Q0R��ZՕ����O�(gEd<*V�&h+xs�>I�y����sZH��a�$ U��a�����P:�g+�{���q���q�M$�F���(��Y|X����>�FK>��\�]��-q>��LxY7b����8�B|�isw:��X|4�xv���P��V��U����t!�/�e� ZQĞBO��B�W��>�Q`_"h_	��E������(ҔJƩO�/�߃�0��:Rq���ݺ�(��ǐ3V��������c��â/����-�4i��v�Lq�0�t�٧���Ye�Q5fD�y#yUHV�{B� ix2�?�Z�q��� ӞD^
u�ү�w�vL�^����}Ɨ�1}i�K�����ߨa���	.Q��֬�����5�1T{	k�*}#���-&�2㞿_�0'����M/�̞�w!�t�V�_��L��J�r<�h�x�}��z:;�ϒ�v������	 ���(���V��X
�	����G���nV4F;d��$�����3u�?�U�Z e�+q��LѶ[1v��ӆUi]
��B "Q���P,�ޮ[]�?A���x��?}�i� `��G���v�\�&w�P,�T���|3KV�-���
��V0V�L@�>�������L�h��w�����n,��h$��*�U��{���*���]�3'���g���p�R�K�`w���ڴb9������,�c����\�ƴ�0���5�����I�7O�˪�A���u�W�X��
�k��&m�ջE_/�a���p`J����x:����S^�2#�J�#�6T�#�P�̲ 1�ﶈ�X���h��U�~k�ȼ�2޲��hi;�b�
H�vR���Sd��r�ҶQ�\
s��36��^񋟫�`K]?��9��v�j�[���a�i�A�,	�Vf�'3�Hg��d����W8G)��[X��F��_^�??��_��n��X7��[�sպw�u�Ib�gI��ӋS�@���vF��7�{�9E~��8Uн���4$e�0rGy-a��~�l���$F�:D�S��^�U�C.�M�Z��\�@����_@!dF.�Y��s�.)[�lA��%�{(�-���ȵ�:�vxtoT����Ě���U�����z��`��T+X+y��Q���w�NZ쇈��m�T��̿�wG}E����z�>:��hĜ[�-�����.�'P䀛K}��\���i:�V�G(�=Vû�zS_�%k��rB��"�.�ڂp��G�|�|��#:m��w�����{P)��S�K�9 �n���=���W@�]J!��w@�����-�����V��L�v~��;+�z�í�M�k�o!<Q�U[E���#�̼�V�bAaXTdR�����]51���?֐ۓ����w��p��L=���J�)��&0�K�HH4�-��#[+X�� &.�
^��^:�Ӧqw�����%��ۄ�w,8���@�)�m�xo�mk��ܬ6�V�*��~�ز��ۺ��Оanr���=�|�fɸ'9U������������MFr��N��Hk�le��8�)��@�z}o<���®�Ņ�,/�������Ng�c�;��\�o��X�Jl���ļ���i�䈔������-�<�����M����0�{\�~N�_��:~�xa���a���cSY��=�n<�����t�M�6��Z��	S�|t?��L�Y8��_�r��u9���ߪ�1�b�˚3l�v�d���P�Cq���ya�&��p1�i�v��j�ǵ�5�f�$���3 ���Y���V/j�}b�:(l��郸f���DBG�hWB��L�s 2Ah6[(�@X������M6��DD��f|���u{�2��V?�V���t�ɰ�+4�z��?|"�l��n�:c�*�T�N��נ�s��E�p�����D����:E�ƅ�FZ�	�aȶ�$�|L9<�Hm�a��4zL�>@�v-�Uq@?O�u8X|Q�ȵ�
��@�u��#�ٚ���V_m����S��c����M&7�/����&�K���(�`��)���hi�,Z_Q�������+�o.�"9W��	��΄�Nc�tOS����^�IY�|��~~^�Q�� �/��bp�L��X��J��5J/LrLb�)k�עk��Ob�-��8��H��X�R>=;�O��Tc�������)��>�<����Q*�.��/�f/mݼ�Z�)� ��Y؟��E��^�֩/g�Bs��I_ݱc+��C�C�e���u���ݷ�6.qzu��n�~ ������Gv��E�q���f�6K���Lt�r��La��	^���������{���ooig����s]�;(���DevĹ.����ߥ�T�ϰo��}6����� Rr�UAC5�4������8,�!T����`؁[r�hԭ�!4�s���-
�D�j�B��1eQ[3���]���8�$��
'��m�l�l:�1<�*����3��V�&cBØݷ��U���T$e�JA��9��'r&R��'+Ӻ�5#m�������k�\}Vj����ɢo޸U��Ԙ�)��p�.ȓ"�J?@�.���(3~_B�����`�U0���q�c���/��)���y���#2C�x�Ɋ���
eJ|����ϛ�ܤ��B�t��|sڇ'Ioe�s<V	��Z�ܢ���d��ٺ +*��b��&�6_ʑ���hB��G���K��N+ H:6,��
��V�Rp���@R�]a g�'(E�&Y'�M5�?�G9�п�ŏ2IR���d��Yio2&l�(f�a^}�dOgևp���dZ'=�|�T�R ra��}Ch~���)�n���:��m��#*E���M;��3M�r�����1햗��/[�`�z�N��������Ȭ�!-�b��`���"Mt�L�|͵����m�sS��O�*AR�yG� W��ErS;Y��}�K�`$�8o/ƴ����(X<ţ�	�w�ׄ�w>�C{_�]�1t1c�g�[�C�XG"��E7���,
���=I�T�FA^�S����}H����/��#�����7���h��yEq^��迢�|�/�Xk,�q�xF���dk/3m�k��V¹��bK^X'������@9͵�z����E;�)R���Zە�Jki��b�Y�Ku�ە�7����d��D��s�)���Fl��I�= ��L�6Χ�OӖ~󑦏e���j��?�7a$�m��A]%�@�@�~p8��a�Љ�kf1O�u�A.�#�����i���J2�q�۱�J�z�ew����#����M�����n&G�"6�"�ޞ�R�=`/�Eˆ�[��1�bx�k������H���)��Oy��~�!-�ݪ	(� ��>�֡������V Y��:w�?%+�n�֝^B����=�a ?��%�]�h��E�"�99��1�h2�iʉi�>�*Ԅ�������]��!�@UN�ŪbI ���ở[�.���ƽ3�����P�Z��?����R�M����/,A[�S���=��g�4J�kF���rP��/�����>� �Nl{wtYGI;�S����Q)�C��e�)Q�U���&�.��`�J�R�H�6�g�>��e�
�Y
�6N#/��5�BWz�J�M��We#�b&�w��J��{�����E�R��?����h�V�qQj,y��`�3	���8���${�2���2��Wc_
lKx%b����.vҌ��7�qdt�eZ��
�B(���":�cb*�#�e�T�;	��8�% _}�|�d>x�zp.��&b"o��J=]w���1���(��p��x�;`��Y���NF������&?3b,[[UN����z�R<e�e �k���ԲCer�&�'׸DZ�;���)(�1�{�f�E��k��፡�������i�6�8��͠����k��B�d�x�AM����d��U]��0OI֊N�w�G)��M��,�>7����S��	_�3�˫�N�x����ܤX�C=����J�ۅ=����H�y��`�Ԙm FI�3�\�Z'1/���LȊE�o�Pe:����m,�/�� �f�'쵒j"!� _}x�^y�?����>�R�)�����mQ���g��]�Sm�zTeʟx�����7����7*:���|���Fw�W�5�n9b��4�IF;��V�^��H��)��Pg�������2S`5��Pp�Vm^�a&�}�V{���F0��������_�;h�hI@�%q0��bmUy���#�����4+����Fo� �Z��؂�P��%��z��{�(�(��N�4�C�Ӄ<��ə��ĥ�}���s�F�������-��pyp.>��T3��_9���'Ŀ��w�����f�
�ӃA#D�+�k�Zz�_���`o�K6��AՆ�~u'���{|O$�eh�by}6�q����X��$h� �>��Վ`�)�I�j�j��rRݣ�s�t1��+���eߓ`B��C��"�,	%��0��0	$�qxF���_�ڨ���?�����^�DH\!�W�ת�&�MG�$y������y������G`�܈�]ș��=��J^p��Bt
���^|�E�;} ����^:`�G�eY��`%���7�7]~-�����H��֊�y����B���M��O��*� ���#,���#tx�͵�:F�.�c����1$�=�s`���UOߌ|�1Ы<~{�&[Ҭ%��g�2�:U)<5)@��A��\W�HQah����b:bÁ04���ȟ?Jк��ʹ��v̇�PE-�0�r�3w�c�Β��zG�|�շ��A�覎H�;��;קr��>��p(�r>=Ż,�' (��2l0%0f�t_�����U�L���V�ϊC�Rr���c��dm��Uy~��M�ճ�E���3 [�r8�w�>�Nq>�eH^o_���N;��w����g��/��D�"�fL5v0�忕�&b�*�M1Aw��e��on��?So���Q�T���.�B���/��X̑�O�T�2i�,w��_	�SD�d��| `�w=��WDd��o��.e`�?0:g��L�zIJ�|�'�Ag����*w����`�����/:st��8�u@�J:��C
�P�I�	��4��KXz�P��¾�֡*Q!��/Q�4J�L��5. ��䱣%�?�B�F���tsN����	��Y{���y���P�6��s���8�qe�a0 ,x��veK�a���p}�!�(7�?�����K��,V{��\��b�~2�H֟��,�{F���x�����W���d�M2Ϡd�j$��'ڕ�?Ps�EX��Ȧeɱ5r���tl`���[8��Z!eN�u��'�e����_����b�s�c����!�������,a;��y=~��5�=��� Y��C�d�2H�CH�,�~Ѽ�S�\jjt�2�Z�J�wy���N���]��qv�*Z\߾Q��X���C᭶�	�8�]��t��/���UxD(���[庍 q����;����-,��x��K��z�59�c���B�����8),N�x|��a�/����er�*g���!�cL'��µ�~�0NHL����5���s(��V���7@�n�Fׄ������(`5R�`�0n�������lab�nG*�>���㭱qk�Qu�,i���F���~Pަ�)T��m��.4�O�7ݡ7�?��$�p?$�M�L��\R�kð�~m}tʷ�5P��<ǐWb��8��K4w�:� ;x��
x	�XW����A^�$�yb�-Q99��?#�\��?x�!����|�vP�Z� K`��u`#u �|D+F~���R1M�=^>nq�.�H��L� �A����!�� ��t	��L�,�;C���J�D$>{����n�~�E6B�!���b��� $�[���*f�u��J�
�!�d�rn���o��x<ѳ�0��`�������Z{
��qFR�&�����V�0|p��B�!�\�P.=7RE2Z2� b��h/���SJ6���j�;��A@�=�P��F�0���r����n�B�n�D>�!���4�F�7��t��*��?���IA@|���;K_ϛ�#|��l�@l�e��ojz$�[�|/����0��\r�bc4rr�_��b4�+*/t[�W���iL�`��۠�8jg�-ލ���:�u)��5�K�;̂����u����b�8�����Q��Q�Qa�����v�)������D�s�J-�����]
�'�I�*#K܀r�<���	�@R_k�uv��ǘGx�W*d�F3���uF��`J�Ø���D^`���1�kS]��"��c�h<�>[��Jq.'�`�A�	]�&ą��4Np9&��H�Տ1��#0�m��y1�� �̡EW�]:��Z_�q�7����E �f+A�Į��)��Ƒ�1˯.�AgZ[<+vf³S90��',5�f�fB�1������������3>�	����ߩ�l�9������D>��3r~���Ew��*Z�R�.����nſ秚�A+q���}��>/@'�tҰGA�!`���jP$;I�P'�8��kɻl�a\�@�ڥT����x�Ϊ)n�XuFu��)��%KE�l���<9@��T��s8��;��d3�၍g:}Q"qt�v6�h���y�NpY�i]��T��۔�3����j��K���kU�%�QȺt?'�4Ր���qW��h-����(�yN��E}3�G��| G�.
��Nؠ�v^��O������TW�����|-pH���'S�EQ�O�?��5�^�� C��6�Ej�t񍃒����w5RB�F{C����X=Ʌ����J�m8EpvQC��J�=�� �\��Ӻ����ި%��\0��/Nu���[^�X!I�婾�lN�Z/e�~<��^��M�����~2�V������G{kW���	�*�u����l���b�4�t�i�"�2�T ��>�^L?OyF���������Y� ?0eu��z��ۻ��.��u"]��=�s�{[�ܒ���85�R5�G�@=&w��T�Yk�B1r;��̪�t�dW�~���� ՟6P�{tJ1�Q���۬�Q>e���o��MB��r�dG[�A�A�EPȏ���~ʻ>��GJ��x�b�#�����5|[ȥ�0�,�Hk
�
z�qCϞ���Q���b>$�M.�/$�y�W�%j~ʪ�����R�qp�v�
�a�U�ò*�ĉv !��L������2��ԀU�v�����m�w�*����S�@}u��]����6�P��g�v�]����&����Tj�(?t$v�׻�֢t���7�W�����i�������[J��؁�_�w_f<�>|��Wk�y�@%�p�EPB�X�ٍ�uD�ܺ�L8����f��ώK��2�tAfs)sV�~�8s�Y���6!�Jŉ� m/e������ه~���9�p�kS�fe���i��D_LY����f��ʑ�*Jآ�V�Ϥt����pɲDL��P�8�P}���l�	�=��;��[0��ӝ��<�Ӈ>�c�`'oO�L#o�1��RZFL&�O;�{;;�9St�|���%Y[FbW��УU��$�H�G%�$@q��<oK������hE�(CW�1�s��f�������t���'��������Y"��n�[��=w�xVaʻb&ߋ��m�"X���F�hإ�bf���1ĺ��_yM�+�%}ߨQ�	?ړ�������@f�Zs*�H9����6�dCŞj��eXfx�UyBF��[j)�oJ|f*���Ԥ��ϮUɍ��ĲV�k9�C4˾��,z`�s&W@��,|�])`7�c���-���5����w��2�]=䡤�_�����w��������7R:!󻳓��Kk�5�Վ�݂2���Ӓ^?C�jtqWCT����?ʿeq'���ǥ�K=��n���[���ɳ��@�$Q���6 ��`}��:6��8?����mP�E����b��E�>f�DH�o'_���R�K�3k+����d݆&|E��_LyWF��[�^�k�Y`��!�D9q�����H��r��#�'��0��y�_�ɼV��A�@Y�������o��W�w�g��p�9{8��)锡I�|@��.o0L��S0�a[ù�?�>�� ��s}��𫷬��䮄�'c���k�K{��պ��	�Z�������i��Fr�}�� :�����&�]�x �$���\���.'<�es����i��ݵ���!_��I)��&`{N{xxx�OO� ����"m�1>r�y����ӯ���7I��0�"�b�4�ћW%P��z�"�<=�T<�?��a�Y\�to����/�����Zʺ��WU�&��4�B�;`���HH�L�*��	��ܹ�C����YX��`l��l#j��ոd�m�i��dsu���)Տz-��j:W��d\�u5r��y��Dn C����3�T)�XX��Ô�����	5����� �Q8@��2o��j����gّ�c�
��\��V���,]S��A̾`�P��B]�^b0��W��X\}��¦<��W�����FH#ە�n�q����Q�U# y�5��*�I�6D���A�æ�`��VQ����U����:��s�����
TVFs���S�]4h"%I�����0�Eª�����P@0^�2�LD:v�]6+�啙��Ӓy�_aR�g�)�g\��>>fڳ]O��H��jqu���բ2���+rXb]�E���0R��B��2��ø�)t6C����i�(�\}]w�Qd x�$A�qL���@݋�GQ�T[1��ol%*�|��x}|��%_�@��АQ,�a�2�R��L�v��T���#N�k?&P(����m�g�YF�-%�h} a�E�9C�ȳ�T�&J&�M��M�H�ˆ+O�/�[c�:IW?��y5�D�/�ہ	�����ϱ���Wi]��
m
��G�1D������˂w��yj��bi>�XO�%Q����쮜�x��S�M.��O-���a"#7����� ȭ6�r[z���!a��x<�*�b��޾����Lux�=rҡ����X�� f�k�~R?�|��	��H|�g��8V����s�}��@5�HEMe����jX&p�*ZU�������P��7�����&b�l��W�Zd��P��䭠���:�
��ֹE��[�m!�N��N���5,���ɼ����v�D����*��W3�9O\;f�C���6��F��k���i��r��6�k���\���u5�|zA�#7Ԍ'%�N�
��E�_dV��&pn`\;�.���&��]I�䌗Q�[����n������������M�6�3J��
k�{Kw�Y�>&�IT�|,��^��S��Uv��5����"��g��g��ao��$v@U:�A2��<�-a�;f��o&P�E�[�Z?�9:��ڗ�����G��J,���{�Q�w�G�fq�L��BW7���q�r� �m� �@���G��V-�/s�4Ⱦ`6�h���1�=��
{"�&6�t_�9��	��W��wW�v͂�;�-Օ!*p�QC~����'�Dv6{��W��-Xu(oc|wDhΨcF6������k��\|�7�{�ّ-�7B���4ϖ��a��3��H����}=M�R���xD����|h���רښ!.%n&#�gCcty"���g�m�,�:��3��S�����ì2���r����`۠�X)o?�c۲��A�d�9������&���G܈��pJtXܐxύ+���� �=9�
5큫�0����v�8܇S?�h��K���=�&��'�1]O)��x�z],����qdpAXK�6����}Bm
3���`��1l.!��9�!LG�Fİ���F���7�D�~#i�����E���:��r���U��9��o�ɓB!�
���3�u�2U���=:ȼ��d�T�;C8Q�F��Mq9F)z�Ëg�m��p�de"��u$>}":����>\�[�0d9�0�C��wx���^yX���&Ȗ��r��v\�q�<��,���"�H
��yH<�`�M:�#���n�/mw��w��K�>�"�B�c�"��V�FU��7@/�_x���h�d����,y
���רe�s�T�[+b�����
���X��+wߤ6;|E}�~[�+8�X���ar7���<�)���ˌ�lo�.7@�����s��z�>�=s�
��/ȯ�%`�#��5K:�(v�ΏN��;�5-rR!�O�j��P�=ԫ��kg���ڒ���H��G*r�@d�������m�@ M��J�ͩ���j���|hb�ஒ�t��<�n,�5�x�n�b����8n�+S܈VM�`���������u��Eʖ�	v�K����* 2��u��ކ��h������KR��d��w�5�k�<]����aF0�F` N96���
�d�t����.��~WC�r}=���r�#n���-���$O^�]�/&S��A��[�}6�%��E���+f9�x��9*�&"U��v��a�.p9�<ð41%���#T�X�1�l�?��WvWH@���J��y�j��}K3����
�=���_�F	x��@�Cd㟃k�<�iI�ѓ'�̗9��v3|��R�VL�T�Ə��k~�؆U�GN�G_������.�"ۈ��gس��e`dZ�B��o�`t9rA&�<� t.f�����	�D������~���{�(�t�('uM⬛������X��4xO�W�YGi��ĭ�e�"H`G�$UZV�!h)%��|��4�ٝƍw�!��%O=�rL� �73{Ub:��Ɣ;Bp�5��ZV�#���&j�;�E�!ʹv���2z�]�N9Ʌ���`И��i�9MB3�}C"[�3w@�0�m7�=�7���}��eYqlh��<�˧j�t�8	���ɫWfg뎼��W���ِ��ZO~]3t��W�r��������V�9����6����_R ���{��Ri��
�ARi
�Μ8y�3$�uB����z�&�p�JiIC�E�A+*�s��j���J�'�E	�R-��O��h[5y���qK!<$A�Tf�L���آ3�� ��c0%0;����La��X���F���O��T�r��;�L:|&B}x(�7����y�ÿ��\j��ͶPS�A�'�  ����<�к[����;P�Q��vٞZ|y�1eE{��Z����X�S���Jƶ}�V*��`�R�ބ*�ҷ��fg�uָX����TM[��%خ�ۯ9�[F#��Xd@+��=���n�$@�/']7Qߤ���hہs��dg)�W��Oo�Ϻ��ۈLB藪�@��nH����sj�u��	꽥>b�=qf���������rʌ �9�F�_ˏ�gsʶ�S*g�ؑ�w�^��u9��`�Y¶�'Mk��Y@>�!ee-�	�M�J����m��x�Ԉڜ�8�m����B�Z�݋�,����Q�4{�m����5=�Y�w��*Ă�$�{(*�7�}���ͨ<�.��Pdc��s� Q�/���I�ٙ�L l���_� N'w��D@Y?n��ʩ	��z��ؐs�$g�uV �ʬ�S��D��;��C�6r�5�C
����aŢ8�Zư@~3�v>u�P$���u? ,*y<%�"m�w0|@��R�2�n�*%`�q?w����)c�#{͠��3�3P��R�T��R�Z%�V:�P)�lѧ���r�}$pr�@�f�¥�QD���s�8��w����{��Q� 
��l���­i�#�2��F� w����_fmڅH�^�G�Y����]�)�&%�F�)���Hj�.���]���[��Le�U	�o�U�M��ub}E{z�'s���E�{d���t��,�Vk��n=kX=Үě@��B�M�]4!��XR'yj�n��[(�Rj�#t(��p��[�����ZD�=(��#��4���t����0�����o��V�U.gg��"�g��Hf#w|������#Dw�%z>1c�MIL/�O�&�^��8����,�l�Vl���#fd��B߆���=�82i �o?3}?Gx7�o[P����:��T?��h�!���*� ?luu���;��۱�;v�nC	�993n�����?�ZRWWB�=H�aw�˓<-`	렝�d��%v���݊O�8uIm�|6S�Z�ܷ��Y^'f?�&��Fq�����;Ö,5:�1m�<�g��[���Pq��ܽ��e���$���Ij���V���HT��Aa��J�~�	W���lɍ��)�q�;H�����1��ڎ�Y?�clen9ܚa���)�sn���#_�/-m�3lVg�$RQ"����:�b_� �榀�Ƹ�Qg�G+!�:�u�D���p�{����|���~��H����cS̭k��������?��ovݷگ�jK��r)ٷ�����|���WIV��,�[C�J��������Z
4���'�"-ֈ��e��T�g�4�R�����iHxV�}�Rh��e�zK�JC{EI׉P�����ccI�@B��T�z�G�� ���RڭS��"��>�^�f�
�&��v����=ۣJ��a�r�5��Q6 P����`�����C_ȴ;m%fJ��e&�J�����|rz��10�m���s󃭽�v���ڟ�o!s2c���2!Q����s�9���wu��sHY����A�f��L�π�OFmwۉ��ٔ����hL.�f�.�M�U�j���� {g6hM3��G�O7[[��>���P�E�	CI��Q�N�GĢ��	USU�o�q��s� �y�� ����:�\�����6,QT� ����w4D�>��5���zy��8���illi՚���}���?�������_��0�I-��uI����w=�����ZSP8��"�3ù@3���C�������-�R"�W?J+5c�g�As�����L���������>�4����X��b�|���@MJg��������I���pb_��j3���`���Ƹ�ͲT�������7��Rf�̳-��&�[�`OgU0�1!���sM<jV�<��w���1��R�Qt)�`�s�<��ِa�Ch#�\&\=�t�%�~�MR�|��f%Ĵ��'ґ�d��c!�o�a?L kn���5B�0�SＮ���Gi��`5�>�x�uYZ��VleP����Pfy�r����j����~{�1��W��>�]>�܃�D'іh����?�4�b�Cn�L��v7�]���m�8��m�~Y�o�as�7^�	`� Ao_����G��c�$?b�#$S�UL#׶vuB2�^��
#[h��9��%�F�C������Ft{���h�Nsӯ��V!A�	^轻r�Pr���h(Ԯ�V��,N�Z�h.9�zt�C(����
U0� �ػ<������uݏef͈Ų]Q�͉!��f�C{�MRT��s[x���aF9��TPn���Ã-�g�H���<���^θ�^������*/i�B}�>\�%��(4�rp'G��,&Y:T����j�<�Q�JÂ�2�F�,�F��'���м��^��t���2)��#��6k�x�tW12s�����:��y� ?,Зn��K,�w
�`N��a⿾�c�XQ2^����8@+F]��U�����ih�?P���3��o���"ˤD������Pz��^���}GIݰ7��9���\�~��fI�ͨ�)�G�RP��Pl{�fNJJ	���)##t~�4m{N����+�KΨ����s��'eSL�j���~�1�Y�q���p�`� ���������o4�]��)���אVABi��O�M�9U~�ը|��T��u���嚦�
&V�SҎ����fc�:r��д�Qy�� ���?�!8��"��&<��O>��F����lJA�=ft9�3�e���"a$=*�V1,�6��@�s�:�n��`x	�6ç��y�)y��7+ra��v�K��-�Z��l\2̦�3��4Ӄ��7�ݬ9����і�i�o1�>�I�x$C�JJ8r��8)֘S�|��3�
���m�x�>7�Z�=�-�ͽ�t@k�+@SK��f#F}��;`����_ $�k3�`�<�Ac���r�8���n p�0~�5����/��L��e�qX�m��bjuu��c��A\�_#S�l��.[F��yAU��N�쿅H���y�`Ko|Z���%=��L�F�L{�wW�~���H��%v����i�<�u��E�B��_4�1Ån]B:�¢�ٳy͕[�G���w�Jh_�t/��d�~�K�������Ҟ���'��yP������v�Lv��k2U�sɁ�{�r�\+�Ոo�|�	�����
���q��&oR.Z֝3����Q�x�(��R4A?��
�]���Q�~�<VdC���ȟ���3���;ME���
�^�q�a|l�ϙ��O�S��Z�d��=`�ટ�sr��oן�⺗n^e�`K�X2*q{�8j�%d�4�3�{��y�y:�g�펀�4�ǔp��I�1�ު�Ɗ���349�~.���ަ^o4��0f�ٚ�\��>U�[�l����SE��#4�1��4%p�p��w�7�.���AKD(�Ɩ1���Y�x#�Y��
Q?��v��!9>�t��0�ڂM�Cr,�˵U�]�/����*��iJ4�R� +�@�)H���q��(tFsMs�=v����U3��?O��i���
�G��7����ŵ������m�����1�u���K�������������������@5��F�͗X�}�BJa�)(U�w�TTM��X�R	�J$E,�p���:FS�I)��[�w|�C�]�Ʈ-r���A-�	�q�9[��@2�_���!�	� �!��ֺ��2fr\��[�ʈeS�m��۔~V����J�7>%� ���+���V|F���9�'�j��tA��0�+zj�I��R������3�)��ʞu�Y²P��\�����*�Fݹ�T�A$C�A'\547n12-S�\��E�6j���/�����������dq�utM�w^"���f�d�)�8gw�h3@����Yz��zW�eASe�:��~���U�6��4��1���L���m��ᵍy ��N�
|g��1N��Г9����vMM���#�)����d|x�&��:st(�C��T�T�,<�u����!(�Z�݉&�M����=Yji�r̞�}���^1�u�+j�[�V�T�I`�>�Nf��`%K	Y���<����;�����P��^w��wׂe�܅�7̳8}�#��5 zsa���*@��;��~dR��UC!�v�58����9���A.����FˠN.��3�X>�����5A`��j�E�Q�p/�_�Au����R� ��B-o�Q�ùC�4�C��c�}	�v7]>�:-���tqqX+ꏵi��FE�o!��>�/V���hTQ/"⤂,� {������Nb5?���_�=�_�}GQ���4i����.9��q����ݎM`agrf����h�wբUǚYʨ���1��6�a�љ�C��p��>F'reGO�v�5{��,�g1~ȝ�P���t�mOQ>��	,_��� �ż�&�8t>IC��7���eH����ޥ�S�S��{��s�������T �M���}�r���Ak�[돖"༺5�6�c��C�X�Ep����˙ݸR�\P����l��w,�c��Ufh�C�^�%pl��Pl�Aɚ�K\ǅ	���c���bU=�� �?�95}Jz��}�&ډ��>j��=�ӿo���kOYj�9Fyc�B?��/w�/��~Ӡ���ūi�?J�}�k�4�,0X��%Cn\�N�v��Q�p���}P�v�����c�l�Pgu�����
�Wq.Eg�i���DF�%���C>O��]�m��OtuϨ�}[qv����'K.aJB1�}���?۞�v|�i
��?64�
�����٤��)�ۚ�\�|���!^�Fg�Wk�8a�h3�T^�&^&%G���-����~т��ik�6Ў"#@z8�	;컋�|'� cpO)��=ӡx�|R����K�)�oV���G�48��8e@��>;q$�"zq\�(���ބ=؃�ǣj�o�_o$���1�|&C�p�Q���'�5<u��G��^Ӭ,%+�#����s�9��}z�����0�h%J���;̚�/��
!�'-)�%U�/�,��6�Ƴ��F!z��DY�,I�n�t��".��0Ȕ�4޽�{�l�%���D�w���Lj2c� aw���+��I��¤q.���J�9D��R*	�A��^rS�C�
��ٔ���x����ɀ�'c��J�]X�X˪>�9�Cbo�`QC�X8�J���ڟv)EuLb5".vŌ�t����=:���@��AHJ[�����]��Hͳ ku�b�	?5M�kU�Dc7���������e6WsD���v?+/1[�
�M�*��x��
F�i��V�ꨅN��zog�i"w~ݗ����g�ʞ��V�$=km�����2�tWV���Qx�DXd��t�1��:�iSG��?�E���&����%r�+!��oŮ�++�=��2�)|�~��,�(�R��~�����1���b�t�P�=��k�t2;헅���RMI4ѢR��_+���ˮ��,�k�~ZB�Z��rB��Ϡ�yi&;9$�Ý@=#��fޒ�ǝo@5��tuvHq����m��hz��v��sc-2TBúƜ�N�su��i
}�0�Ap�|;77���cL� �s���YR�������z�`1��;��s�Fw�u
=��DmJ����_C����.��01A��d�T/��rW���+������0�ʊ��{�� ��JU"Wo�,7s�CrzJ����;��|+R����io�Dz��{�aM3�e�Z,�T�,(�v�7�6�y��1��s�E@�D���˩�̈�G3�@�J,d�T������J$�^o�Y�ʶ����3D<h1�Y�{���<��0}��%q�L^����L�Q��i��{�s���+�����+E��{O�(@"�ƀ�~F�<꘿mA��O��t�g�b��6�Jl�J���'E<�H�|����b<�	W��alp$�7<�
D���u�ۙҶ�������;7S�e�������`CMt>����Q 1��#���r����A���a�hLZ{�5dg�ɲ�cI����vZ\US�CΦ{�1��HQs=)K�Cc�-/��)��P��\�+o2��Kٕ��;�VSov��A��`4��B1j�9q54%�pЁX��ڎ%ۼ�ߺ ��^��	9�T�w@ �3[ݤ(n���ܳ��70���s�p�
:�CO&���<pm)�*Aq�ē	�A��LA�ϛ-�>�f9�5�|���g|�bTe��� ��*�Ji�з��8�`�Wb��"���G,���B;��O_�=7��צ�BM��iuǩ����O�߁��\iq�4w��TO�-��Nz,��-�Z��)��g꧖#��?��\�xT3���5�y�?�$>�g���J��p��P��T�Uժz�9�mFO俘�� 'M
����Vmeyk��0f�`]f�׶Lr��}m:�yO����EH����R0n��j1R��ժR����i��ݘ�r=K���O� *Z}]�ߙI$�>��[�C�Ï�D}}G'FMU���񓥰 J�1����9du�_d��������8�̵c��p��2�O@�es�M�{��j�>��ʯ��O�vRw���
�R<���9�:m�1r�~�ƴ0���r��HV/�N�dEV'^(��2"^�a��!��'z$&7���`�N U�gh��K�bU���L�vAg�+�p6���'w�W�$��HU_���~	j�C��&�l��c���wK��US����xwQD��fi�.5	�ӝ��;��8E�[R�F�3�� �5��<� �������H����3'�k��z(>�F��+�;8n��^8�/�T�mN���/x�J���5�:�w�S��/Éx��L5�  �p�X��V� ��j����?����GHE5�B��
ΊPT����{2�]�x!����|�B�Ǳ�@��@
�D�u(#0�a2��,�C9�+�a-x���O<�*��T�w��'<����Bl9�;T���]�����y�%��3��fr����8�� �IZ&Z>T�G�8�\5_���?���W|BJ�%ZċQo����A9�}��V~mGO��J�.�k�
��=|�ޡۼWmqS�j�h�8~�ҍ�̙~�s1Dh��~0�*T�Yjƛu��AN٧����ӈ��޸�&t'�I+��L���u��qiȮMYw��uA�x���r=�,�m�Z�)=��,E�;a�(I��h��PS{X����v�t)�9n,퍹��t7.���FJS�(��Z����a�\�Y35	A����J�:�7��nc�n�j6��!�b����Ot�+��`D
�5��2��">;�4q�# 6�f(�nw���E�b��^������,k:�7-���ހq�D�l�_��0�_�r�9 �>k��(b�	>:c)��i�ꝈUU�t�B[����Z��m�.���,w ��d$c�J�#Z��A͞5�=y��.ؿrG�N�(�m.��B��7j���M�"S�l�Ȼ���xΡX>3��� _Q�b��F�%��{eX��[�`����s��z?��y�&���ޘ�t�0�S䳁�.�����c�w���%7��u�c� R\+�1�|C����@��ʂ㑞�8m�-:�/�kmᇻWT|��i9m�"������%�.o;Sf�T�Vs��0�j��G�P'(L�iE y=,� ��	Č�p~� cC�>{T/s�/������9��:lt;�۱C���,�M�L<�����oC᠐
܏,s�����E"%D���Vg>���G������o�B+�5����ܶYj� q�)5�d�܁d�Z�#>u ��*�2�k���F���0%n���oh�]�uJ��!6���j��4���>�m��#��R3�}(F���.��k���IRs&������
�X:� !2W.�ƈ�u����`|7e��Ҍ�Ra�HmI�k���I�P����`H|�sw�].m0�Arph[ЋFТ:�D{���51�j=��{��(��+����1ت�֋�� (��$F쵼K���m	�C����{1'V�(����1K�/���^n��1FߵMx�޺����N������_�Zy?T��Y�<�������4F�L�"�˳vvrq�f�`���A��Z��7�L���}�b�!'���5Uon�	l�s�(�
�8c�e�3�PD���M5ߥ�釂�M��PO��]��Ǝ�k��d�1�O<t}�2����.VM��$�`%;v�A�$�����E>C�)�=^B���Ⱥ���"[%;��'��x�����q|�& -M������϶.O8J�B�>������*-��FK�=7�p]����-M> )BNga����b��M� ��=Ћ��^��&�lEd$��f��X�v��0��N��^��Tb*�Q pC�Xb����Рt�����N
՟�e�I�.��#��l�����d͹��đ���bk��ڲ��%���$�h���"}�F#^^���bIe��|�l7�����gE�(�QM �8�����*�Ǩ��-J,����	����XYy�Q�	�0�@��.Zt�!l�+�7����'nT`��;��"�=��&�� ! Ե�m�ᙘ�r��PT%I�7�J��&*�]��֦To)�K��.	'_��	ie�?�m�?�"���E=]%���l�i��BrR;���
�1}t�&O.g�XHk`YQ�[Xi�Y�d~� >ۂ��Ӡ���]ȵGK3ǓG���w�QD��7
�Ɠ�-JG�Ж�j���s���;��$���Ȩ(�~և��c��^˃�4��ܗVʓY�=f��S2έ��-�+ޘk��ڼ�495q`A{C_fR/����3��!(�T�)�ӣ<m�<�d�@�4�H@�ᦊ����wajN�� p��0� �@c�?�b�gQ�]I���U3路�>�<���D���6���0� �C����m?K�I�<�V�V���~��������#� ���J�V�"��VԈUd�s���4��|���ы�����~9�����`���S�7hYC�!��@ٻ�U���d�����	��?T@��Q�g��aa�_.X��J٦ƌ�����r��̞�f��-�#��N���E;KR�eZP�g_��Vu4,l/:Ѷ$� �~�1ϵ;a�x��Y�`yB������p�mΘ�d�|'�6��'�6��QtHb-�+}i�y�P�e���J�-G�9D���D�P�ӛy�y��Ѣ�LV#}�W�7�aH�G��g��E�*�m�%�!ξ?��Hno@�݉*�qOv���>�v��?�U6�Mn�h�)��Ge�£�<��

v��~�G��=~��j����&P&|�m�w�bͦ_�m�er>�����y��*�ǒ�[�G��{�~��/��fL	9I؏��>uJ�>YaFw�R�#=.Ѳ�W&p�	�\�
@cl;�8����9W�K�h�g�ӷ�	 ~�Th�KDwh�� �z��2����1�K��m6;�A����A*�2��6��̒�-
��7�!�z�����5tN�*�R�n��<���ٷ�|8�:˕��F�A�j-܀��Q��U9�j~�{�td�͆�.��i�(`��ĺ*pV-���\��OR���O�i��S�C�����+��.���$�fP5�p01��?�d�,�L$����p]x_Y�\.}����6������wD0���U?��|4ڍ&��$������ܝ���<��Q����Y	�0�)��dzO��lSS$(Sb�Q����Db�֖��V;�5�	p���q�g�.�w�%=kT~GF&N16���Z����my*�A6Xƪ���YV�x���n��&o���H#G����Ak�����u���J-1t���;|4�z1��������(��l���V���f[�:P�D�~y�^QN\������m���?A#��%�K�곉
�Q�@Ҝnq:GK���PS���j�z,_IUBل��&��Ƥ�����E�?���f�-4{��H�x}.����� |Q[O��V���-N�J��qt>��-$ľ�o�:�P"�K+8���u�����Q�:�e�-{x"�N��#d�s��G�������vi��q�	�j�<��"l`O���5Rƌ���5ft�1��ެ�Q}�߹��O*�����	���=�Ǭ�<���/Ѫ1DP=�$�&���g	�.��7"=�i� �ӿ���dwP��
{��a7��=XJ��6ӥ0O��4�#C��1S'�(9��]�n
R�G�(��^������̋�� 4B[*,N�c�V#� ao��B�g=�I�},����܅����+e�[L��3�����1tꎋV�N\)b�XP��^��L]���J�<�s�AY�Pc�b��ff��n�˾R$�J�I�W�2��萏��3$p�Yss0m�
����1��7@�_�煆�}��ߓ��&gy�"SY�|�z�A����Se^�Y��(I��ʧ�I����w�(ȵK-�g� �x��gΐ*���xz�?�X#�ֳ�� �~2���%\+�{d��v�<;�	U�N��<{�A�ਙ��*�[9�|�m��P��$�I�f�?�	~\��@�"Ut���[k��!���x���p�� BV�hc@ �Y`Q�`w$����F���m7Q��[�`mt<���2�O9��(qi�yn�������z��H�x���+���1-�S�ۺ��w. �ᔈ����9�z"��եj0?�{��:�
W#]��f�ìS��,�r�k|�zqU�RU��q��9�u���.�fyB8�Axs�	�q1Ŗ�~Vk�y,��m9���ۦ�/\�Iýi��o�WZY
zK�l�`�PE��\J�/�$ߢ�������)4���~{���c��</�2k&�|P�bh�*[����:�\-,,�^|����}"�vlB�/�U��dF�;텛6z����7��75K�#�L�!�ıx�����^xb�Y���^�vj�'蓝��;�B��b���¹`>S�ƅn�����&���&�/�ֻ�V4�'g֪��z%�Osb��G�>#M~�*"Z�Āa��B.1Ͷ�:O�Ȁv���|���>�>����E��zSx���6���� ��o-�#��C�ғ�1���1Vs~V�.!�+ؗ4_�̎� �dN����ey�&Y�m�ˬ��*z���y�o?�n�po~�gx��^�sGj`��'����8�$*@�UhM}�_/����8k5!�br4�-cEY�#A؆��T��Ѝ�1m�_r�Z:�(W�����pɶ����(�	4��`�0i���U����ע@�%Qfp�@b'�tX���������J�]663���ځ��\v�gv��z����=��t������>)xж��qd6���1#z� HIjz�3da����+��
$�I1f-�H�?',��94��r�%[�W��β0�r���9�^9|z�H�5T�Cjy���1��j7���yPFZ��zp�h�:_�I~鷕_��:[�ٷ�D<	�]e3^��0�e�zGy1�Z!H�J4�v9J���]z��|G��(N��Kf~a���ܴ6��:hq���>_?�q,���㯔��{���gƍo���F?���`����G�2\g�����a�.3y�Wp<>v�LJ�E�C�������{��i�����h�)J��d��������c�f���& @L��@�o�Q�������B�H���;�Z���,�1�[	�	�hW���T��ݍ�U����O�^��A��wt���q�]��k��V��Ī�s������5.�^Qp ir�Z2jJ8cee��n4�ڽ���8��gf�eW�#�c��:Yx1.g���O�`�w��N#������f����|vn�lw��I��˼�߾��N�{zu�^��2I\6+�QM�G�Z���lN�����c�"�W&>N�=��ҧ\gj�S`�T�h?_t�J�,�D�!k����S����8��5rA���'Sj�P�]��������)8[G>���6�P�ӑ}�1^8۾l��{�?�	�6��d��U�=�O0�-��_�B��p�p�\&B�bg}��w��9�2Z��[��d�4]�aE�.���ܓ=G<^�a�Ԑ���ݱ�N!h�w]F��dS� �� N(�>I_k˄7�կ4��:S@A�VB��f�*�U��><O.TV)N��wpl�xAHt�BO��U�h��3oY'�{#ھv0d�g�Z�FC�N��$�uWD�Z��2�q9?u�xƞ0+�k�b��3�v��BM�L[��*|�x�j�1�����dC��I+�b �1X9�t���yt�����__�8���%K1�A~*rH��|1|�hc�_��W�P����Ea��2y�l���ZMKG,u���A��y�C�V]���r��m�7�?���kβN�ed����d����B����``�ո�ز��E|��%�:�~�����̍�5!�HF��2��2���QM��M,[@��ZT\�͉���s����=�O�ْfDȊ�(�U*���5l�� �k��e�{a�q H(kz�'>0�	Z#����V��O#g�$R�,Zv�M�'�\N�y	h��EH3�8c�!��m��xD1�|�������0$��T���I*?����#��W�u^"�6����Z��ü�NG*�b�"�ߧ�kA���Z�$5�ϟܑրy�ެ����FK*��Ui�AKR/���:E�Im��޶�է��d�#-�n��k��]�7�?�NAv�1�8�e��ؽ�?�� ��؁���GɎ��Ɍ E�ef<�fc�eo:=��V�����Ӹ}��[�t�W뎼�����:���P���l�k:R��>B�.Y'Ԥ�sk��r�B (S楚)l�Y;�?\-����J����YT< YՏ��AR��{����n0�i(�G�9���c��H��H�`X X�D [���d,�Zw�)s�ѓv�4�6Q xĕ����:���`�u��!������ ����R�f�ў����1�J�~�5��fs��6A�`���j�!�fò�$��LN6[wQ�����~���֡�R�F��T*F:YgM�.�JZ]�����ά�XӜ>��4�ȾQp%!��`F��xvOv���W��f��+BG2�s͞Ő�t�m�Y0}"�m��x��a�����z����.�k�Q���'��@�db���Jd�WcOj#k��јרƶ��C~�[@���k$�WHE-���[����bwn�k��l/<6%�&7��.���ڢ���OP*�޶����W��~�0f�4p�39so��ޠ�:��fo� (�4�Kl��U���>U#�m�^w�SƑ�2g �3\wC2�ͽ�#x�g����
jo�ğ5�w���,����:�^z
_��FV(��47��/~E�tUۣ{��H�O�z	�/��u���4��U�G��ŧ�g	���.��<�������D�!Ln���$�0P&���Ӽ�E�Yp��N��%	[⯪a�_����
��p㷱�w�+^㢗 ��>wHx������C�P=[I����kG�rn����
LyW]�$�%R��5���2��.�BMɶ�6YZ�	�f�J�Փ���R�^��:�{�f�����ֻ���7������ޏlDP-���l�3�>���9.z���tF}ɋ���W(3����h2l���*`��S�]���L
���I�2ɕ�;�,�Y6VI=p�̮��9����T�=��N͡�  [	p-�4��\��Id|FV�����C������W� p�H��VmL��mجbn0�uՑ����D�_K��0�NVr�6�ۏ���Y`a�����Tmp�]���tZF���G.���InB/a���E�y(�dr��=tNw+gu�6��?|$�2�M�����΍��x�Ǿ��1�$�1�.�C��Q7�N7u�\&O�J���%��������!.��p2�^�@�b8Ju�f��q�Q�#�AнnޮƳz�'�%�=-�Z���D@��	�Fuw��C�~~�6��^��(�������bbss�l�G�P��e6J5�����Ӝ�$R^ٙ}YQ�j�[�I� �ft�9G�OvI���)Q�����3�=����clbM��d㪎�s}ȡ���:�n4�K߲7��2�(�/o.�d�F����h�������'۪�4܆�������id�"�ϺF��&�׎/Ė��
BfՌ�
S��P�;�)NX�U��ǵ;Tvq�������B�;doZ����º?F$�v������A�ٟ�Iߟ,��9�:F
?���J-���ы?;��|����F����|�������놣�L��_u}Aӂ0J�	*#}39G�8�ɹ�h?�a(ߖ}��*5�KE*gauj�W,7\�>��t?X�?�߾��F��q~��i��a�Ω,kr~�ټ=��4� ����|5�z��M��vC��*GZfM�?�p��x�O_KQj�_]�NX������R_�]����L`xwx��Y MǍy�c�CJ���鍮�@��Kɋ�
���Pc1h�Y{}�̢�M��÷�ѝ�]����MG��W��Sfͱ�|mE1����큇�CUv���n�)�}F��S,�L��]bR�Z��L(�)W�n�\хbS���D�7�VT �����&	2w���$� ������d����p`�>�uO��a?߲��׍�I��RKP6� ��.e�~���0 Q��������"�_����=���^Ͽ���@��s�]����ɲK9}���g$�f�۳��7�6���I\>����*�5"���p	_�>���mȔp����Ӱ,�B��#���.�-0��YL{�k2�ĝH[��&� ����-Es|�G~b�Yg䵞��r< `�^�),w�m3������ٚ�q:t�ȹEx�W�t�Qɹ�+-��D)uo�2���7��aq�g3�ޔwYq��2��y��5~J
��#��yX���!�/��Z0=#��ذ$vGR�"}��N�쾈���5#�y�j�N��0�z{	l��&�DOO�M�i�5�l�|���܏_%o�¾˴e7L`������k���m����r���|4"�e4N�eT�6M'p�7��J�=���g/���لx�C�N.����<b���kg����ڀ�u?����}����7x_��������6�|nmD���ZϬf�'g���M8x��4�:b���~_Α�f������~�O�)�����Zr�m|��_f�e�Gt��꣎Q��b7Cf�����6��ȅgau�+�/�\�u�x�`Y��wa��!�{t3МN��	L.�"�;�%�跹[��X:���4F��xd��9B�ɮ�ȒJh�1����V��X�:Y�i2G`�ބ2�"���W���ٵ-��@��=T5�HR�{
��-�,/�)�6�������l��-�X*�QP�\��ގtKP�,mSp�'�� ӳ4��Vt�6�"PpF7�����}�a6:��0��S�+�5�׭yM�[<��=� �@��mHJ|���7&3^���K��F��cW�����Y��\���i*�A� 
;��M�Y�\S��
��e�,�p�$z���߬��462)ݦ8�O��T� `��&]rN�#������
FQ���vy>Xz hY�KD�z�,h+>�N5�NyW[�/W`�q�Y@4�q�X���L�t�yw�\�sE�N�+3�+2��!'gs���\����w4�Σ����A���ן�������B:Oi���J����R�1�F�ONgU�Vi��tµ�
���w�����H��r�T$ԦIC�|e��,��͎Y�G�(����X��R�(�������p��Pa3��x�����W���w�-�j�&j��ڿ����Nk�6&F���j��	Nv�	NDvz���Nl��x�J� �}��Q��n!28��F�^iEQ�o�W��P�1�?�pj���3������%�-�>=P5|i��D�o6�	�imqB� x+6��R6{�M+�z3r��0Ʉ���D�H���ν�kg���d���`��L�0_ÿ�K�r�b���:�M�beP>.��V�0WU9D���abW� ����̹L�)��h}$&�8f����u �S|��U`#�?��@ǰ�6T9>y�}K��,,d����2H�b����\ts��_w�$��\��w�6�œbz�s ���Wk�˥��	D4g�_fg���ôf�xQ�"�ɼl���ٍ��1a0�Os"`H|0�����h��|��\mKV��B�
?�8nU����A����szB��Iy?~�'�^��>ۨ�rh�%�[f�;�T����2����[T�8�Z�\X����rIA�j�1�Љ��<���_�MYjuz&�٧]� �&��w�x5�~�[�S��~��A��i\!��'�[
��}�rHgiB�oO��`�eSـB�{���t\����I���k4(�p���mN3���3��Jե��G�Āk�(���,�U[���|��6n'������Ɣ�ۻ�0RmZ�il�k<��:7�"5S���B�IQa�G����a�,�Y�)6
�1$!�����0^�@�Q������6b�-{,^�FD̤J�؉�똂��s5�㦀tޝ�ѿ��{�w��S�ڷMJ��ퟓI������C��o^3b޾[���hλ�� �=����T�:h����'7��4�\��O�x�o~��9������~⫦�I���X_��^_"/�>�d���z�6���Zb�[t���t� �~8{y�.O��G[��X��C��`�ڐ(�wj5QE]Nz.s�1E�=��Oj�-��5���ez5j~���@ۂr�F�!�#H�h�/M�L�P��\�X�����B�TcN��v�6OM����v��otS���x�v���[���(F�ݹ�u	?γ�mHB���.jϚ�:���r]>���@�44\�5E��T�d!}��[��b8�[O�+=��\�h��8�t�=ǔ�QD̘2r��0>�@#��C�2XVZ��JQ�p@`�iEՉ�D͑mT��mh��ˍJ�.Y�^h�^�g�
�n�Fb��C컿�7���K��%x�	U�������ࣖ���]+8!�M݇�Tm^W6�y���#��Gt~	/)oẄ�iе�^H[�!���<��Mݩ�N<�<��P�ܙ�W�Q��1�0ݖ˦�D�<m#�`��a"�l#.@Z��6�g��A��j
⏃���ݧ��l��p�У�uP�"Q �K����'�
�;�}H/�ߐ|=�{���^}�[�-�L.1mg��}�чUn#�EB�D�g��27�eʉ��,q51��g�P���-�����^_�=0���}I"#�������c���%n�o���uf���)	2b"���F.A�gM���Պ���Ot|ʔ�D~v)=U�R��́�n�Ǝة�l����B]�NOL�O��d?���7�?��%ꅟz&��l�z0wg6�U?؜�̠`8w4w�4t�U^�^���$t�z��=@���"���ֳJSD"g�|�]�I�oT`��7��)B��'���E6-R~�����+H~�y�3eXE���4�'�b��ɰ��(pw|�4��nb;:^��O�U9�M!ln9� ��2�m��do{�\�C�c�&�[����z{�r�}V�g�ɷ�)�N-T���vo�W�%i{�����������TiӐ�5�I��t��䭓����($��(�-/�{���r�}�Hv2�L��3��Q�̸������K�d�|��irF;I_�.o�9��M��;�;�R͑\Oϫ�X��H{H����_�=�2�ޣ2�!�%�E6�Eֳ��T<{�4�?d�?AݼU	���hA��k���cN?S�ؤ5�nb�����\-���H�a�����5��Ŧh ��Wh ���ИA2���e*�pJ��XV�����L^��K]9N{���ǰ_Iˈײ5�_�e��2
`8N����bπ�� �4{�pE_���YN�(��)|;]o�ʲ�"�-6�6��1��Drn��_�$%Q=�b�`<�$�ju��2[�f�F811�P���E�&#ZTE�.�r�H��V�Fa�6��_wg��c�Zh�����T�&�+�j��'2 Pz[����x��Y29sZ��#zf�ܛЄ�̵t��E5ȴ��p,�?Y_x�l�BJ��ѡ���;�;HeL�H�ux�Vo�~[3RMN���\�k���I�Fdn�d��-������A��&��Д����gv���E���><h`؁�=���y���[��)��R��z\qV��~��ɏ#�V{�7�B���/�@�x�I<�Ə��vקm�#.��"�n��g�bġ�����д�U! nr�.|�iza�QzG��b�< �$	߉�P�����a��b=����jY�G�$�M�U������� �<����] &��C��wY��p���5EI����wm�^��d�b�m��誴�_���\���fʡn�^����V�]�	Dm�I�rb��mXv��pq���@�"L���p��C�Q'�m���uLp� C��ӫ."��p��S�J���z��[����(�>�E��I/��b6fn�`�Y��	���9�YT�ϸʞS۱f]�[:T�4��t�R��06R�k��>!^�T<��ʌ��Z(ݶ��Ԥad�'������i�h�e�`�5������t�q2����c�r��K7�����JĨ�j�>������z~]Zw]}Ў״��	�{��zU, ~`W�:�=�=�u"��b�)��М �G�b�[�s����P��0��C��te�T�k/=��P����B/ȣ�F�
�3bu�� �ԇ��D
�
O1?���936*�{�r�4b0�9���Y�̩:�C5�}#��،��y�)�'$�w�-��[[�{�oC�oc�9iǱ��������U0SՈ�"�Dz
�}iw��Q���͓ *^�:��g��Dx�����p�^;K��)��n�I��S�g��;�=
��sq�
�](�!���q�]�y.��-����m�?c3!��)48���(8��B'�>�D����~yp�����R�U�C~g�M��Q�0P�����u�SNVB���h��iksl2읋$o����?�\�5����N���Ѣ���N�^l5�q'-+�G8b�)���@�@G�)�S#�C;`J��d�ʾ�
a�hgf�J'b��ޟ9}��g���$�Ո�b�[a��Ac��r�o�ŀ�"��OcM��W�h$þ�E7�p���Ic���U�ͩ E�Ρ1��'�q}l���� �I��f�qB���#��',�������VV?�}�E`�!8
����A�:/@�BFR�©gɑSn5h�ƂOh8�6��&�3nd~���4�<�ܰ�p���q�B��4I�b���ܝ
@�����H�����~
+�	u��21���鉿�+���V�{�5�0���,�Qi2�9��|TPb?�g��I�`zs�H_ʂ=���<yz�"�7Z��3��� K��+|ǹ��g1�;�04�DbE6Q����X�-v���SU\�Q�*��	ơb�\���Gc<b��t.y��y�p�tȁ���ű"�y̑~\�@�:�oI�����"@Oc��O��'�q�>+����gԎ?c��ߘ\rNiji�����&�����ܑ�+=�'LG��w�0S,-n�w@�� �c�Z���Z\�_|Do���͕V6|�!ClI��{B�v�w4�h��,�2�K�Ьrfs�%�rx���MΗэi�,�_�.��iu`atI������L�:����1^:/dKR�f}���V����H��'��o�}<t���
���M)w��*bL	���5���e�݅c�v�+��/o�3��?����ֱcc�b���3��jk���OW2�3k�n��U)��t���±�:��0O��m-N��-,2$��_�`]}���p(G�Yȕ��?1^���6��m?�<�&���;G	�%�CZ؆֗��W$���(���8��ة%.�Xw��b�*Z$��ɣ*�F�B]?l�H4'��<S��?�h��
�lT�LQ-�����F�1ɾm�ւX�MH"�{O;�jP
V�%�J��0B�Cݸ]j�者����r����G �!H~�6��s��YT��qa���"TP	��[m>������Bu�x�E3U)��JǗ@m�G���q��0oE�צ��lW"���XԂ{�t�F^7 �i�hP�P21r=��L�D��aQ�;PJ5I-uO�������q�{F��-a�<ҩ������$cR��Rro�TQ�>S]��.�W���0���I������v��yٵ/�P�ُ����R��0��*9�$��?���Ϣ�
&�������ӌ�^67�"`BJm �	���^Qe!n��ܖ�Ŋ�>bGvӱ��m�D�&R��B<�f�����5�7"*�k~�5U�h��G'�n��?�6(�a���j��X�s�,#��O9�2M�š7��+��d���p��:�Dt<%�#��������w��1�#t�A��h���oۂ�g2o.�Q�2��O�誊��k�ѱ���u�k%jh�]�v���$�g�ۊ/:ڶa?Ɛ|vH�~��X��H������Lp��;�'%���L�c&g�-_J�b��_�b.��?�&q(s3�0Žu� |�̦9>�,\l�D���(j-���T4�>4��=�yvXʞLz�~4�s)ae2>�d����pߘ���g�h���q'#wlI�q&����>b��f+W0�z�Ƴ+C�����e���;D+�_�@�~Wc����Jۦ���gЄ�L�j�lD*�A�8j���LOt�f���/I�U�N�TY4���6�;h`&��e}�����̨}%Xp�7���&���������� �!�Ł�TP�&X`7��C���&�Q���t����PZ��@�MY^�Q�����u��m���_ �� ����β$�BA�����vd&�.����������J�Ԍ��h5��,.��D�_�V��&���C	�hzG��1ߛ�V-�����K��ݑo{$��$O)��}��@��d�z�	�Y��	�oݠ�o�$�����	e3�]�cU�R���t�q��V1\��UU�yP�nk��"����W6˵���X�q.�R�Wp� ������p��8�)&f�#����ܠs�3�N�����y�������N�_���"���p�,K��b:q��-)�4T������:S)[sOrgɳ�ՁfW���/$���%�9<�f;�/�=|�*ك��C�g:�� ˭���6�U��R9f�\�s�:�d�(�+���n7+�.��'�3f}{���
ݠ�O��[�Z��&�@�{،�! u��ē��[�0���*�b%�cs��B�p!��g�h�Dp7`ٳR��\01��v��9U��^F��u�KGW��C��k�*��K��Y����7�wC��͖�����iC7�O���$�����7�e"-dx��ƍ�!Y��fr��� "�X��>,�����y�����U�{���,�p���&��i�}����g[�T�JL\��+��V_��4,�`)4�x8�Ȯ�~���/N*�7{=C�����|��[^�R�>�b�XFa�2b	��SS�[-��7��(b^W5[�YMK��h1�*@v�5-o��ي�=�z�շ/��׿A���/��<;&��RŻ��8�2J�i	��.E5Xlz����_S���]��0^	�Y���˷��¦
��t�l�z�!��B
r��h(J�c������o�r����f���c7R��- ����I՗x86�X=f-�~��8���Hg�	�L�w�N�Q���"cսUnA�,����֕,/����$<�LvL�1	z��d��a�4E�9b7?r�CМM���3%�*������Da�╩�x�L����x�<��ҳ�=����ڼ@6l��&���`�6[w���i����I6�+��(�d��+dC��0���9jy�b�Qi��G8��bP��R�CK��j]T����ڎ��\
L�`,�`�{j�7���ʹ]��IȘ(�?��b.�ս J���ɝ�f2���Z1gY{���-�h&v�x�S-ao�&W1{��4��y{�\�����7�^h�
��uo�(w�;>|}`��{� �a6�+e���Q��g��k�E��z����x���2�u���f@��?�Iʎ/���P�9@-�9K��'0E���2�����Yt�șELR��s�}E��­U��ٲ�Y+�駉�:�ܒÇ-�K�ut}���0w���_�iQ�`Q0��۹�{;�ZaGi�y&y���9Lŧ`%W���`Qu�bir�;.��"��?�@=���50^�H .�5���]����Λ�����\��H��~T��.9�=)b����p6k��?�nKg��5��>y�����@��4Hཥ���w-�9�dtУ4��S��:?>�t͈Z[c����xyL��1�A65��ou�������x�I�_3�8�j�n�,��w��������R!Є%J���Ne�c}�-�(���ȥpM���%[	f*#�{%r^��S}) T�i�x=�ss��M>w�5�?j����n�^^�A�7蚹0��xкNx��0�i�i��G�/ޚ���6%����l�;�$)���<H\P�
�3�W���_52�5sl���+v(yM��|"Vq/a�x
��)R��(OS<���3�[�O6@o�;�%0�A��C@ @I1��I0�L�F�-a�A��R�
4'0��F�������0	�q`T��&5��N�K�!~�'����vARt��:<u%�B�_��D�E��iX&��L0\9s��lx)�L�{(�l���^u����U7�����i�oQZ46�f"Ő�4�X�e|+��A9�W��e~���t:�)����=���+	�����X4�W�����t4o��1O>�iӞ�߳�Z��l9�4!Qz���X�
f��O�ai�*]���1_�6�����5r�m`�?��̰��Pr�����,�ޭ�J����7���� ����}�M��[����������`��@l��E��y���zgb,�'nr#@�~��4[M{�pY;��jÉ�.�d��-�6*���2)�J2�볯�;$�y'7��]�g�:oPiλ��PV�Y6�s��b�LkA��� �X�w4���)�wg�]f�����`M�UVm�D�C �`
q!�JO��x�^����e�*;}<ź$�s����v:�2��}��LL�;�D�Ȗh2����qE�ED'�G�����&�G>�]ӄ�_�<ZZ���G8�׆8�4�﫧>�yK�2��;dmG�N���y��"��)����e3KG�"��U*Fe���X`׸�@��w�fQ?����^�L�#������>����5�Xo��̧ȅ��u�>m�K:��_a��_�e\�-�ʻMo	�I�:Z�f�-��Ftk�B��>��w�؈����g��2a�fгp�q9�L��'ּ�C�e>m�m�a"���NH���j��;-o�Y��U6�]"����2���ÂC�J�L���
3W�H�
���<B$����ƺ�
j�'l�֝!�&>�p�q>���)0�(��n�����$��S�U}��,�C�y��{�Z�����$m#O9��*&�U;ڄY�8�I|�����`:��|��l!O;��)�E��7I�^F��a,�D)1���y��F=��^�X�Q&8;�W����������'[���D�
X�R�����,�T��2[�,E����S��6��yL$wO_i`ZJf�X���*"lN�=��ծz-������n�$�n�2m�?Ksԟ��N-m��T��W\��~�_'�,eP���2��� �n�<�(��}M���$����{:���v��A}،�3��R������(����eE4���/H#ɡ"��D����Z�)�͗�+I&n�i��������*TAs�*Y��1��~8��e��l�lYd�|���Ke�]��K��QE�?��R.�E�$�^������oA��[M�35a6E��K�3s�A'a�b�#D96����]��B��'����I�Sjn@o���1��E̮�8t��&$��$$1���50���Io�D��TB����V1�=����������aBY���O�֪4`M^�lUZ���q(þ�
4Įt�ӂ|O�5�fҞ�jJ�l���;�>n$xB�v��N׌���$�/-!/2��z��l����W^D��������2�
�B3��S!�6"�?�3��g�-��>"�M��f;��3s��n�:�_s^�\���b�����ڤ�GVm��}��r��
���Niɋ�#�E�z�א��,�3nQ+��A��z���e�08��S�Y���a��I�*)�b\�.JxwU:�A?\�Xx��l(Z����`�,hbsm���3�L�MP����]3m[H�45�f�a�+rn>&%PJ :�����X�:,�=��xw�Cj��J�/���!�0Wj:�R}hH��_����4���tp�b��#-�4�[Vu]�˞D�Ny�ErI��|�b�C� /�tN�Yq��{C�G?�5�3(��W[��g�C�R�$���a'p�|+$�/!�����v�e>_���۠
�d誮%�[/��e�5U�b��Z�?0�a��}�HZ=D�6�K>:����jX�)\�Ӓ�bhuW��Ҭfc�%pa�.�aD��xf��k�bu�ɼh:(�(W��*��I�)L/�x��=���¥G���RX�ly�6�ɉ�cW+UZ� ��)j�젭Q����Ǘ�m�u+$
������&�(�z�?a��I�!~�����k����+ǳOCQ?�Ub)�X5��h
�ý�}"��OG��9E�����	Z���i�G~v#�N�eQ��E\匥�$<}t�zu/�<�����x�C�����Ef�B*�%���\'�mL'���0R���L���̍YX������)���9ތ�j5�����>E��(O6�w�� �ަ˧pO2�,w�p����b�d���)�/4!/U�+�+����݊zX\�l��%4	�
�;��m��Y�&;'i������^��?Pj�0Z��Vz������g,&�s�=	�kl3�<ܑ� ��l\�2�hGr]��!V�`���N54Lls_�D(0�6ye0�t����@Ps�ƛY��?W&� Z�כ��B���l{�#$�.���l�m�eUEj���L]�_�� �	�e�+����S�0�m]�'g���-S�!��J�hx3���[4���*�	�C�"�`>Ϝ&����Q�«�n�2��@M��&'
"
�5`��ݷ4���z�c��}^(����ryԦ/�z9!��+\�.+�'�A�R���.A��lnǽ����ʇ�ʌ�d}�����C�Y-}��(G\1s^��N��������g�����P[S����h���7�^���m@ٸ�,��r)�R��Xl�qf�fV)gT$�l�+�V��3+]֔�����>k+3K,-E���f*/�.6F��'~hԺ{$W�/x����Z`�^"8�c�vLP��vq1�\�=߂ .����ϦC�~�H���K~Cن�qt��U��E�3y��;N�\'�	2k����D5�=�$g��M�d�<��1�T��^��l�Z���dd_].�R٣|��&��o1yԨ�x����\5[����f��xD;K�"�����ٱ�Y��_d�����B̀)�	Ԗ�M���a�-e�	�7ڂ�sc���kI.A *\�'�U	`gd�<Sd��%_��e#ζ܇�M!��]�X\�ui&��v`%�Ԅ�!���U�Jf���=�����x!q��iiojSXn}��Z���qq�w��p���ŏ�.K,F��<D�����Q�&R�
���:��+rg�z�ɺ$�Ǆ3Fw)�QF��Dd]��i�Y��Ǯ�`�ѻ��f"���Ms�|w��1k�����)_��&����>�%��=��v��K��f���&r�*��>o����]p�+.$S��1ׂ�m��@�+�"��H���7�A�Y	P��aȚII1�'�dðN�+��H̚��ȸE,|��%�R\��8�= ElY�Ŋ!��UE�}I��4଀; gN�u��P ��^p�����3�}7��������H���?��cW����MX��ߜ\eK�_��e~o;�N��� '4�pX��3^�p�e��+k/�%Dl�7�U��T�%��6x¸~��r�����ɵ?"��E���H��E(�}~?t���b�<��'4C��zh�l�M�P�#��q�KVa�TX�{�z�ʹ-�We+x���P@	����M:� �;kgR�1.D��y��*�����A���#�!���}�NԨ�����x�%"��S)����򿠓1���CPn���(*�`��?֟����w'��8!pC�H�7����7����d�/ mI�^g#�?���q2��+k��Y::I���i�=n�����MjR-?劻�t.Fa���`0賈hI\$/2`#�K#Ё�>�+�w���;f\rs�9�ϐ��z"i#��g�V����_�4�d	����Ƞ������֫9�#���\��ǔ�7�%��`9aEd}��-�Ts=���T��E�����֭�,���Ć�	�7X��ԗ`a~״#F8�y�j�CnJw) =a�F�!�E3�2�)Xɇ�s�$e�
����`ԯ�J.���|[u�I�q�sW��YQ��b���y�N��;��ڐֈ>��JE!����l�:zp�VW���V3�U�,��50��v)+�����a��a�RX��z$�[������È|E��Ĩ�|�N�'��dV�:�dt y�Y�}��CH��q�,-2'�Z����x�T��5��5Q���=�6�<֣��K��wi����w��ltA0ဂF�D�\Y��цy����0��,6E���)���QU!v��i��פ[�F�]Xz�t��<�^��w?�B82S�ϡ�/�j���/���I�|�8�"�V�1��n�͋7�2�d/���+C�2��f����I�Z�H�Ts
l���$���p*E�9�%N as�i��u<�SަF��4p�{gщ���O��,%�����C�m�U��iX2�ֽh��#�8�_���[`�.����lQ	��y8U�[m�\��Nj��.G���<'5�o��c�;
Z�S�c�cѥ�4�aK(TC�%c�N�)I!�A��^�?�z�[ʇ{_k���!@L��G�G�"G1.��<y�����
%���\=����m��������1d���^��K��� �P����z�d�� �����ǁ�̝�)ԍEb�k�K<�d�Dl�8\����<�@�N5nE�C�m�B_Q#�` �J.B��+/��{��lnk�^fl��6X8�Ζ���Wb,�9�"x 9 n9���t:- �NLЉ؛���q�a�Ł7B*��ʬ,��tY��=H+ �,U��P�^G�0�м%�	��`\Ǖ;��k'3�t�fKq2c���J�w�S+D��^Z�<����`t���a���!�oCGg8�b�H$����2�#�n�iv���
�
Þë���������F����Ԉ�fZ�c6*����N����m{	!�h����O���x�[8�u|w��X�M#\Ew>�Mp���it6�:K�o�{$;���־�a�Js�vŷ��������b��	���[��)Ư�m��\�ߔ��[4�vtU�G�WmY�@�F{#&�"����b�Į1�7�Eݱ�e���^��$�A����F|Ǘxg�l�p�%?�E^�ˊ�ٿ�B������f?��4}�T�N������Q��@�=ud���@w��E��bԼaW�����O�`����n�]R��I��2��d�Mv�~Ǔ�ܖq�m�f�9k;ܔV�SܨK"�s����VjD-�@��:���������`6�3RU��*a�M /<���t��&��|۾��@dZ�:��%���9:϶�� F���;���@�M�\{�b�Z��A�K��!��@�?�SVǼ;~�=���V�i&�Q��,���c����.�`�dE���ԷRu#�շ�3�߆u��x��G�rC��\��T>)IX�|���+l�Q0��*@+����V)�渃�D�+����
�y�Z�S��2i�T� P@3�*k(Zc�| �-_� �9�M��p�����1��Ų�>��\����</�d]+&ZphJ]��^��s䠖h�`ZU�E�o�ݯ3}<H����%9y^f3�f�;���*e�Qɚ��R��ǚ�T�ל�uk�fs�i7͒��Ye;v�!ևq\��-��Y���6M@`�����c]�J3��o�?l�$�!0�Lǧnps�`
��q+~�]��Z̀"U�k`U���fF2S΁����7�u�0�z��';Pհ|m��}��zh�u������.�e`���۬�Θ:o��5WV�h�Z��8Lu����O4��\�f�����D���\�	1��l� e{@����x�Goq������K.�����T�.X��!fV��1�G�W�w�%w*����ê���b������3G�Y��8/�hhd8s�/!{q���_�IYN�jC�s��(p��I��)�}	�*���i9L++ӗV	L�� ��lz�B�kCT���
�=Q1\�	��D
iEO�H^�_�������ko �[U*��/@�/P�"�)����1�g*����!wg�J�KC��~��mJ�[��m�X���>v^��V��ݹ+?���3[@5���2*�QO���
":JGhɥ$\L���� ��@Rd���Y�t��d�v�@(2C���K�v	ը����-�T�K,��	��=�t�m&|��w�4���5�%{�5�i�Ԩ��� ��l���a23䇒w�SwI�)�Df���Z�>�Nx}��F"Q�Vn�d!y�7����%����#ùVJ���x �rb��}�*�|&�7�a#�ai�P��Y�(R�
=��%6��~>U@��\�a`�pU�ú:��-�4�U����Y�@���)9<�--$3�9]���;�J`s5A�/��=�����|y˰�=)!ӗ��F/����ٻ��ّ��O5���Q�&�Ƹ�n�te�o�A2�h&)����|J~ִĲ�d���Yo.��8���1�$q��r/���D�퐣{.�'dQ4���T��9��X�w��ZG��?�5���U����.��s�BHWYu~���`�9�uѣ�9,�~2�=u0B��!g]�w�d;-9̹`�Xj:¼�F)a��<M>����Ԓ5L�V�lq��G��#+�������8�)/�,M:�+��na���(�E�=Ў��`�E"�y��:�O��U���d��$%>�-��#"��n{��2]�$�>�ݒ#Ʊ?,m�#�ëTX�Q<n�Ⱦ͐��q���)���$��F����8�!(^�$�������?)�CX��_`ju�!�ڧ�<�_C;_�fO�iQ�w����q��\�?������M�E^d^��"���\X���s8 ���z[��z�����}�:m-��.Xt�J7]��J��ReX���]�
`@�x���ے~�4mst�D�p��2�����b	��?TA�ה���P�tc�W�UaJ����ԁV�-.͞XU�-��Hg�"Ǟ��	�3���BËcry�7Y�E���G6P&tm��9�=���k?���=���')���K�E��*�JIIIdD"�ٛ?#<XH����@C�����c��=Y,�	Z��X�7^$pO#]�
(�wfnH`�lm��&hp�Y9M,T�qB�U�(k}�K�} �sueBHc[Sn.�}�'���.���Z���P�,�4O ��0�g�Ჴdx�����I��8��Ēs��?	�0&���1�fk}ۮ8���6VD��"��h�G{u��?xә���+j4eÚhX�S��OgJ[ӀRn�>�F�Ew[�r{�!�GY�5x�tXk}���+��TD;�>�:��tj��;Ln���UK/9(�1����I�
.L�ߴ��R�]6�adE6�">!���J���;�Y@��%��yy	¼����!Fw�����~qMg��h�P^���|��ݥ��k���*���E Joc��<��NQ��
�kv�I��J2.�F|��{�lM+�#{���@'��ܱ�h��W��
 �u�y��{|}� ����r��{Z%���{E��6
<_5�\������k�TW1�bݢ\��ً���q��XD�f���CS�K��\�?%cIF|2�Q8�23i=1� �<~�l�j�3̕b�v̂���6����Cu�n�_��v~��1�ej��a��Yhd�ܹ�_�9�=Jѷ�Q�e�?��T�Nk�1��z-��ǣ��%��kW�W�٪_u6�I�t4߶�$"|=�s5R�)kr�K����wc���^-�:�P��� f�g�B���Z>6��ྕ��p���c,��'�a#{�qΈ��%hH�H��*d�^�}1������t�:�r 4,*\�*�s�'���[���B����[�Q�=`��-�~�GN1�yX��z� S=��k�ҢԮ՝�%2I�w�@�,-�v�{v`+>Z�p���"��2�5��]VZ�괡 �T��1�	�/h&{���6�	�U�5�;����ί%hi���;��cr�.��g|����(c�!��GkV�Y�y5�Sj��}�j������?0-��F��*΁�(��J f1��4�],���<�^��FWE*�So�#>��(�I5�Oy��K$��K�/�,�L��+�/��/.��=����s����r^Ҳ<����Ò�����=������qD��9
�.��������m� �&��k�x��������k���7աٳ�\h�І�@�]r���)�+'C�+��I��XnM�G1��Qx5*6�#�//�χ�c�-_cH�sl����oRY��-�T�,��g���-=��n.�S^m]�6F�wG��!�;=��`Ӝӡ�d��Z"���	 Z���7��H�M '��{"��X���s�C%�>�����d��A:�ChDo]i���F;m'�<r�����zO�宋����kOA��䡼y�� ��;p��9?7� Iq�*r>}-==�;<Xb-]_A�|�B�=(��fm�
��҂d߆)�H.��+:��k�N܄w��Mpc�=�t�Y�(z-׽eG�}l��qLs�]
�9>��aK�$af�����y���
��&s�(d:!pY��W8�<�HPs�s��h�m${��E�miߨ��덤�6t��s��(6�Y���^
O�#�B[� ��LsF�P0�_��R<�]�p6N	�ϚmjaC%s��2%M��N����}+4��O7�O��{��Ջ�=koI��[8hW�9�[�@$�tx�4�����B��onH`{*����[֖�b��b�<���I�a�T�<��čo�E�w�τ�ݾ̘����*<ԤgK�QC.��JKRSR�~ә>�4���5�V��5]�փ���W�Wz��7-�O���?Eu�w�N���x����j{��q4%���8�Bk8t�ʤ�l�Mоo3Dz�	k������@:�������PĿ��5�U��T��OC�2n��_��Z�o�X���VN3��qe$dέ uu����X�w_�������e��?���R{�~��ބ0���w�ziIWپ�Pz�ŭ�:qvW���+�%K�ip�=o�e���C��ߤd��y(�AE�+KD1��p�o�n�ӎ�H]Dk�r��MѸ�y�+к�����0<%��U�!��6����+ ��j��0��g�C��O�d��I���.p�;�<K~5Ӟ��}?�y��c�����e��G<�5�ڐE��a0
VJ�k�uV�57��_���'����vJ��R��f�V���F�Ũ9��$]��=�X����u��6)���!�fVp�4�n��T~�Ӣξv�u��1М�ɍ�*�Mw$�3�?-V��������@���D����q򠝛��\�ҌK�Z^��I��aA���@ޱ����ߴin ɂ5ĉ�5i'"�)[����mm��]"˞x������Z���*��<�k�]V���G��w%��!\�~��p��I	�(�q���>��x&�]� a����O�W����b����}*
�]�	���>g��K0�[�`*��q���)4��Brg�涡�=7J���va�f���	�F�+ ���ߧ3M^`z�eQ>�g�n�p9�b��c.�tc�Ѱڠv�6�x�2��x,������!���i�h����`��
��]��W:X !��-uG1f�R2�b*�D@�_��J�էO��_�O����<b[��LǕƓ��)��?.|�k{���<�a����-+̸ta�m��5�u�ڐ��I6��я9.;�>l"�օ��1���D��|z �C���aAaC�n� ������#ˍC�E���;U�h{���+6)hUk���#�r.rM���I���ش�C��uHv�^Z��/Ms�r��2���k�7Di<�}���B_z��=�R	K�z�E���4Y'�K�#�F߭�nľ��ҭ�D֚�9�����(��An������4[s�,ސ� �T��i�|+�_�3�7}+�v�I}�@���((��.�S��Z�@���A����O���D��FO6Pz���V��T��WH�	�+�?�>Yp��e62ƵR����*~����g�0�ڸ~�C�㊡��q��O��K��줲���6n8���[d5�6�}�_qi�6A�/>!;oXG%�Pj���- ��Ǫ�k'Z�n>P���;����96f�6 �o_�F�N��X�k���1�$k��L����ͯ���C�H����+���`�fOVіcOR5"F�����S���T���g5tI-�����LX&������&��Z8(g
�g�E2��ޒӘ��5��o�z�R�оX�
g���U�>'Q�v��OG8��s�1s*Q�'�����Ӥ�ej�߇qik����<Į�������!��rû����~oq�Q2}Vٟ�y,5����	h�@�\��'��.���)m!_q�ݐ��/�8 ���2j�3;;�O���B�0����4�e���n=�֐��jTY�k�H����Q�(v���Wa�p��L�2��aʵ'���K�&w�@�8�U+�Ѧ���Pa�m�"��jI���8}�<5��g��?��f�Z��.���pɸpN{=��`��6L?_�4�3Q�= @�M��` ��b���Ϣ�<�꿶�B{4�R�YN4�EB��H�p�*hV�V;�F͂�2�bZ𚷜ù���:�GQirD��#P��+�׃�N?�gM9���� ��q��PC�Ozuy���U��h$�Vˬ0���+�r�����ӐA$]c	�{��� ��Y�^���m���E�wB
�{�R���j	�_�G)���O�9��%m@Y��a	3���+@�b�\fk�����E����.���FVX�/���ӂ�a�2=a���oV �)�3}!�R~ujB�N2�ӓI6�M�D{��q|LF�'�S{�9�=ؿә�W��іW�]�O��X�&�w�H���;���G�I�A݋U���G�R�qQY�3�����^���-v2q�#�U�2�U�_�C-���N@t.�.Cπ6�}�	�G1w��V�@��sO�j�-QL���"�����/�e�,��3��t"B�os������L���wc���m�:;w[ 
n'���[M[w`���^I�� ��1�J�jq�)��W�Rn�c�i�iǿi7�0�k߯�v��T'���$�|*U��§�?�>�h�������W����&GE_��Gw�%'k� ����`�,��Q1jB�ѭ@s�^�㑘_�@Z�$p�������qC��s��u��'�5�?�v�ݏ��e�f��K!
9�hjp]�Ȋ_Z�V���Js�=@1?њ|tF&v��E0�-'��|��d�@%~`��eY�p���uw���r5z�7�^��@����Y �馮"�{"�i2P_����^(���x�����Ǳg�A��{-s�!����[�'��mE��$5g��;���A�ͷ�1�t�	���.�psϐ�b�i���ߍ�{g��q����/D#��x!Gp*z�e|��:c�1j��&r�Bѯ(����+���I��f6�ۇ��eR\����Ls�y��2�qb�`���E�{v�'p>W4$wXLg�`6�1�@�(��|��w)��9B����PvnL"a���=�шU]�Q�ܴ}��AE�ty���vd���&��Z���(:���q�9l��-M�hO��}�OBfK��t�/�K[��ؓLf�ƻ�w�s'�ocdK Ii��iF�[0TN�����[f+�r��Ù�������2�qT��vY�~�<���N��y��B޵��ȓ���:�[�}n���^Ν�o�#_����n�']皶o!�eu�o�`4[�� _�8TK��[�!
ʌA0�!�?��7�*������)��d���c��ڍ4Py`|D��L�:0L+�z?�>s�ܝyZ~����,���{A|b�Rp-�5l-.�� ��~\���MaJZ�&�7�u#�X�X��!prkIy L]�w�3 ��چ'��K���������@eʌ�������F���xب�����ut��Up� ���b_�e~��T���K��R̂��J���YI/�؄�^P��b�i2�Z��L��UG1�d��r�hO �7���?�`��(�ڔ�*=JO}�,�ڝ�Vu=J�g�f�	�6�!>^(��&J��;E=�fvY��ӒP�O�6�"˥r�iq��-��o��c���ǝy��}<Bd�o����{_����UC���ſ֨�ğ��^���T:�H>�G����O������?�;�����%��'Bz�)�F�>>wj=���ؼ1�[�@.�|5(�>�ԗ���krIi��\,,69���ڏ~�@��2�=2�hT��>�'g�%�:���%��f�������xS�qiSN�^�z� ��WHH£��0N��"�f2�\UCt	ˍ�g
�J4k%pҙ�Ğz�M�S�(�)1Z�5����z��^m�j��[!ՙS�2�i(1	������^w��y�V��3x�j`nȕ{x��%�[��$єH�1	�4�s���{����r(�ZB)hu4nB8K=ofu$���a�UPi��ԓ9��P��w����Q캭J�D���N��l�p��G�kQ�`�ޓ E�*�ѰN4~Cـ
��U$y۾쓜Q]P��Er?)��A�.��c�*z�)s4�LR9���qb���ra��0�ƍ��u�Y3��ɬ�ӛ$\/���f���a�+�֌���(&�,��DF}�G���fV�9K̆Zu���|lS�'�Y.��x��"��U(ux,���l`s�[M�G�D����._�Y.Zrl/���Y�Ǣ��R��:Ke/~�%r�ZF�C��gp=�fՇ�
��Z�o�s�����P��$*m���x�-d=x�V>߉n B���=��x`�Z���w g�@赺`���jTgmX�)�5sC�i-��NlU"�r�g�,��	�.��=��$JID{^�֋�U����#ԉ/�$�iu����c�o�L�,�����٫Ec1�h ��Mq����H'�s���If�v�L.�K���-��օ��z{G鱕�hzgG�Z������͖�MD��U N4�3F���V*��7�s=Ёr7iH��H{H��w�����:i�>�g�n�U]S�T����K��Lpc�ɥ�4
Egh�y���a�����O/IeFa	�qo�����������]|Z|&�U���Hڀ��K�5�h�#�L�0�}w�/�aA��3����1/��Jx��gƱ`�H��H/r�>%�7!8":Z��2���`=���q�ٰ"6�]>����<N\bԻ�\Or�i����'�Y�xItH��A��*���Aoyt��-\�԰J_R�YҺ��x�B���TS��Z'�Ti�Wp�FeCl`��G�Y���RU�l|�"'��D�4�^�zt_��DV���65��{Q&ʵ��+
�+���P>����^ �f{[�UV�lW�Wc�ئ_p�7C�(XV�o�t�͏��i<f�%O��ؼ�9r$�Bh++�H�	ã����\���	D/�V_<ۨ���q�*���
΢%:r�X��F�Y��a�W�B�=�H���&�Tlk�[|S?b%#��O��_�.���"n�y��Y��;��� �y��tQ��{f���l���_ZC�0 �-�RNhK�:��'Q�yl�٧�����ԇ���d����S��'ɺ���j��5L��pH��!չ�e�S}��3���~�A�ls�y���v/��������G[�#�T��-=WБZ�U�l�S4����:qM�����jF{vBl��~l:zA�b����<r��oRAU�D+���p���nq��[k�,v�M�+=
%=M#�|�è����S�&+�tw�z�zTޓ�'����E}��w����s'���#�b�D���)�u�ye�_��B>�D%��Ca�P#�@��cƼ�*DK�- ��3^��i�7�1��z�&e��RK&K|my�k�L���y6��fz�@�*͝å���@d��}��_���M���n󨆦 �*J7��I�An�y��y/u��H��D����W���\���'��h�.JZ2��̘�l2�O§R��3n�`��Ι�ǔ�_�2�j�ť�]�7E"�s��Yյ%�PsN�+"Z����=�;�L���(y���������\�����ι��<���P�,�O��!�)y r����א�9��z0���O����e���7�����轩07���MB~67!�����'MT���J��zT�)��x�K�A�-%�$�DRc*�M#u��=��KF�M}���4���댤�c?}�R�v&B��=�L�Ӳ���d�D֗6�-.]z7Жn)�S,��\&R� ;aRȚ��t��������(؆{��5#+�U8OQq��]u�51�%Ӎts/����qk���h	P��j�%�+�=�7�.���~��}pS�����-�m^al����~�##ҩW�ˋ�lY/k�Q?�1�5��$�\�+�! bL��+|��$$;�ǣCW��_��D=P��H�nЮ�����~8詳�P�X�p��@���.Mu.߻�^�Qމ����)�b*�6���&��5%R����DlȰ�tvs�*AD+tw�+!.'$��Xw����t���k$��L��Z���:?�S�_~A�"x
��\6D�*������NF��O)���{v���h�q�^����-�,tc�gٹ��HSG�����&�`'&�u��޿r�Tw�0mv�Z���%V�z�CO�hG[N�+�p��BU}��T���r$[N�pƥ��&�Y84�����3�� �N��I��V���_)_�,_���N�*+&`*j��%�Ma��ؓ	X�Θ�̪?桳S!�̫�"���K|B�u�AZ;O���ؗ�W0��a�\9�j�-���J$����?u�]�v���Q������`Ƃ��W�U1���=�#��X5�r�5�}�d&n��g��U��׿�<���.$��KT��fhu��_�q����U}���P�m��4@Oc�Mn1')}^�^Qea{(�oR�x��Y���ߩ�g4�?�jm��I�[=��&�;�8[�l���2�Ǭǭ#���7ޥ||C8�0��n���}����ߘ�v+���mۍng=��sJ���]�;�:`�Yg�>'�\�}4�����.Z4Bf *��C+�}�"Jڽ�o��2���Zé:��ε�zO�8^]*����Uw0#�(=p����m�	�S��.��%|k��K	&��pN�����y��xr_�C*lI-�#%}�Z��0���\�Jw(�L�x.%@?�X+��Z�?aFnس��pܡ�F�'����l�7���xrMܗ������@���ɋ=�$H]P���A6�q��d	'M�J6�g�n��!t��M�dW�k��}�,_O'ڪ:YhD�R�E8p��1B��� ��G�8����!��[�]�����C��d�/�AMV,�F6�/��o��֚T`�F�c���v�l�P�p����@��=��	�-#�ߥ��c��lQ���R.��uDV:Ŋ���Dj[�t	Uy����w�#��QD��a��1R=ftv��tP��?b��sk�Q ��g\����O!���Rq]��.���ng6\oх��#A��;�3��Q�J�e�&q]7��\��R�iM��Z��Z�G�<�c���\���r��
�����ɾ��A��a�!,.~ʆ�o�̧0 ���	��tF�}�����/�wx�Է�=���L�ʰΌ�:������ɛ;��((֩��35�'���m�zZ���(��b@�a� ����❆㚨��r�_VQ����c�WxJ��O��7��c$�?Vec��"oh`��m~�!hL-�nR(�ސ�ʢ��7*{���[���8��\1 �7�>�+.jDP�cJs����Gy�Yibb��(ǋv=H�S� �y����z_c]x���\v#-� h��TU�v�gN�\F�7��)��Ty>a�Z���&r�]���o>6y��L��&�s�}D�.�
ouŁ�j	�*�� ����)$..��=��2Ȱ�M���� �r ��� @�%m�"��4��y�(�<s�H�ٚ}A�� ��^��Sd:AV�$���I�kK��ޢ!����a˺Q���A��',���ܬ[�q�n�}�!����z� y� ?\���n88�u�%S�N=
\/?��\0>|_�Ʌ[��;���~��v����(�g��o'���^���`��*^<������#��ʤ���'�c- $���F!��~t�k�����#q�6pć����5Rxr2V\��i��)�j�V���ٗ�ɋ �:n��d�AsL�~!O�|� �������QAw?��2�Pv1R��ii����x����[e'l�zԬ_]󀧽^�:aL/`���^��W�ۍ��c���橰͎�j��X�k���w��Y^K�[�&,Q��	��L2��_VR��Z0
�H�����th;œ�I�/���e[������/�<,����g�k�#L<��o��V��eb6�6��]����r���P^YZ���m��d(
V�r����{Q_����c����M�Xy�v�mh��j/�{j���VE �����
��%�V�u��Iɖ� ��V�;?������� �y[���C�
�s	��	]�X �A�%bc�����fX�u@�M�d��@mƩ����?y6U ����+�օ�Q+
�{� W�.�7@n��|I��}y<����f�=��������F�,
&B�m�Wé,)�� Ft:p���@�P���"��S<�hu=�&q�D��=���Lz@�Y%0�D��
�o�xo答��`eLM-G�� �������Kk��s?��0}8@�����s�^�Y���ds7���Za�^v�}��(�J־�p���!����5�4��P7��**�XoO�iV�x�3�嘴\���i��N$d'��P�Z"�Z"hy�:[p.�aC��j%ѥ0i����s��cd�����V~AaMg�R�R���Q'l�z3��K<��2�(צ�;I�#3]y��f{;>����A��	�ߌ�M$�C�9B���هEɜ��۹�����+e����b7�Z�q�~`q��������t�������Fcb>enV��̟Z~���7ZY�s9�pj�ݪ��w�PxXa�o�$�qvκ_o�hC��-̫衐��K�4���Լv�	�,b��$h�1S;woӟPXX���U�
�di��;Ŀ?���<��4�z��;���A����VZ�� ����N��g{��+�W��'�@*|"�����@��2�o�*�w�eT��/��X?}�`Z}�hE��j.�1b�(I��ج���d�~�^�u�k�%S[����1�Yf���]U$f�m����?��ǅ�A H��#�O�ȣ.�7!�(�tӪ��v���EaL��q��E��1���u��~Q7����M"���b���R�#�̥Om�q���������c��^f�QCi����	߽��,H�*Bg@�����=Y����ے�K�ZR�;c'���Q�D'��٧y��wD9�d��D*-��џ�	��[xM1�91P"���ű^?�X�#����)��IҊ�U\�"40X+���^|���{���?�O�}]��qq.=���#�~�"��i��ܧZ�p3�����$�J#B觪�Kw)���Z:�{!�N{���#x�_4v����4�g8Ə��~�� 2���i�5�mC�������k�H���nfM��S���^ ����o����ӕ�k).@.VQ]Ck\�͢J�l���I���BgZ`�{��홓!��9�i���I�Ѹ'�d�*x��M�=>-�>� �GKn�O��aM�")�#����yH��8�����I�,`�˻	�������,B�ŕp�^6����0�3S��7z��k����-?�Ϟ��ڽ\J�<5.)_���[���օ_��y.R��.k%����sŌ"��=C�Y)V��`<�SqW�(�\�|Ԧ[!E����eY�S�&���|��'͍��c�9)�X�<~��bW�j�lTwW�oZ:�q�3:F7�Vj��x�JY
�[ƅ�6$u�f;J�o7T�ز��ͥ2�Qt N���zR��@{
xlbb�[��~��XMD!�jԦ 5k���I�ؾ�V:=�E#�H@�_����H�C��,���NG��c2E�~q��a��A:��ċ���Vk�NN�Hq��MZç}���!��r��	�^�,�6͚��L��\n���; �{ 7�	���K.P����C����XQ+����H���>F,w�c�{�1?b6�=�j���a�0oT�%BS]o�}�W�Fm(�!�=��iP�.�:��qW%�@N����᾿?Q��IjʘL���Q��͒�Ҍ
1r򝒈7��J���rx�gݖ+6��f4��N����|9�t&iY��j�ӡ,�]���]���,��D���PM��-�팅?s*C%�F�]J��P�\4��4� ���� ��&��l)
�؜�$�b1w���C54�����l� {`�"�U�ZCm����ͣ=`r��x:��O�)�[���6�
}%TWS��2)�k"�$��Y��~[þ�Y�"�{L����a�tG*G���n4x���$��'$�Rm���~~����-#�%mH�u��2���axT����VLTb������Y����/v7���G׀�8Yݎկ~�:ؤp��B���c9����A^P�2_ֻz�}��ܽ\&���iq[sW�<��-P�=�~!^U�V��W�Ƿ*��x$"�$��y����$	:��nk�RԹ#��P��~1���Ouٳ�����ܡ��W�)������5t����c>�Č�5�~����?mF�n��D�o��'�E�%�_i5���:����R�51Y�70�Ǯ�q)��_�0��0wΫ�����yW���eK#9�y�^Ql�e|kh�bl5?f�"���lY�U�G|A믜ZhQ�$�e�;������$�v������m�vK�뙟��0p?����i4��8�$<�II�}��du��&�?�\�c���C��`*Ϭ�?���^��`�?3፹=7fCѶ����L�C`�j�:��.�}��M�r���tB���>�s�H�Q/G���X)�����2�|'�����eZ�S:�U�*�A��Pov��4��%^9�1%�6��tƑ�1���2����w��}gL�y��-]Btl�D'Y�y-4��zt>�tk|�nx�#���X��W�E7YΑ���h�ݪA÷���.8�����Տ���i�xd�ӄ�&��e	��g�Û�� ,��R�1�)�囍�rNt���5���W5c���i?7�&B� ���V J/��>5�4^�p�x_@�N{t�Ʋ�2�	4]/� �lG�K �P2�(��3��8f|�'���#��7�B5�y4�0�&�"w�����\�����blT]��T�>"�|	*&G�S�����|&>��,:$���m�n�O�=3Ը�62�j�(���Չ�U��)�n�i.��tZ)NI�Ҝ˥@�Z?_b����/��k�?d ��k����H���y�!�3g��������e�@�S�����?��d�(�$���FȮ�u�M�	��S�n�Kp�4��R~!��E�qZ
��^�s���I{�m�7�c�7|+8 ~.I��%�i�mYfp���iK�0s X����#����{����Z��H��3�S���FK;��<��'7��n!�x�}�`o����V�Ǹ"p���ͺ��uu���`���B<�����@��\A�`�{Gk�O���i��6��W�#M?�#ֺvb���;܋mj���NK�N!7�7��̑d�ٔ+c[i��AH�%6��x��^+�v���~�F�Ā�0�f�X/�Lb�p7��#�W�U��0P�'�.�8zmx��=�`"�JZ�w�Sj)�F�߲/~��-3G�i
P8��f��i��zq>y4'r,f��?���H+� A�_39��1��c��3��xrl�3`�-�zZF���)
�wFN����3D��:�>�"S����I�yD�`���;K��}f�Ã�C�	�?����G�r�s(-~���F���S�K�߰�.Z	딯�[�o���9*��ٱD��_�͂N@�= N,h��ժ��rt�Ɠo�m�cͰ<!AX[p;��2'VhG9<���C�X�e�E��B�_�>�܁�x�"�����RUH��J������+����6��O_9�b�e��b`�m!�mH;a`�W��5�2���toak��$�Dc`�JW�]�"~^���7;�$�l�k�J���V�n��#ҵV�HI��m=L�*ٓ�������`�l=��l�,"\�A�kS:5�1�ë���[!ڲw��98�.j�O���n�^j�nK�������6E��}Pa�0��c ��E�O %�6�]�7d�|��R�7�٨��G:�K�R��ά����|��}:�en}8�wP`7#.h��;m�`�"Eo��nׯ�aP=�4����rh��R��ߴ�m#�)��O���/�RK��C�G��뺍�� HO@�����ʊ���2�C:��z��߫��,$��
���4�漠��[��\�%�c<�3ը�?�����f�S�q|ɴ��/|ui{�t���)����ض����͸w�\�t�Q��JٮwY���QGtqh�~�D��8D.��ܼwnWpwRN��f���Sd`���������38{�N�[�ւ�sk���ط$~_����҈�b�od��L�9pO'ri�-lX<B��W3pRo1?����c*eM8-�<�|��R��#�!�a��?�1'܌*��*�9��1&�9�G8�jx�J��˝�����WAMZ���D˗ ��q�����	9O-��׏�2����j��??�ߧ8��U
���G��'�O����8���]��--��w��;���Aj�!D�MB�FՋ�ٗ��YP��j���patg�a
U <���/mZ�M��3������7e4h%&,����\�!Uz�քG���C��;��/��C��Vc
]�^ܧ��%��!�~��k����kj*0���]��fNp�a����%�(Šo��0cH�F�. ��	��/}��pk�7FEOn���a�3���v�5 件�w��4�����O�rUN��}������u�  f
�.��2$�zh_o�n_�zA���"�ʤM�B:L*����%���N�,)g����o�@:|�NY�$NR�f��Q�y��:��i���)K3�0#؀�%0�@X�@���iE�H;O���9�Z�u"�� |`0H��o�)g��@�f:�{�܂��J��V������C�+G��Fv��bO��u`)Y9��M-�p�[���mL𿬯n!��~4�k��I�����dSG����V4t��X.������3U1�B��#wX�h8���>�>���~�ɢ�O���G�-��iJ���e�������~�V������YP���*�9�y*}}��y��j~OC�%�*�������`[�������+�.��v�����{��5HwP�m9!l��/7�f#��ܦ�����R&�E,�J}1�b�ʭ3�}�8m�(>��Qsqu�d@B�ꨞ�̒���[Z���qh����-'Z%��>ȃ"c�\��)Y�?���s�v���}2nl����dO)��|S�W��_���B��lc_�8�2��H��q+Io\��}Q�a�~ڎ�E�V�=�u��B���uLdK�C�˽��Ȼ
9x#�%F)���nP��d����>@�w�\��@)�Z�� E�@��z�(Ҭ�C\���ʎ[�+�=	�)����-��D��~z#:����螎v�/��tR���EXa^��΢��NֈFQ<�� z��O*�*�D��<��]�>�
�����\��J��y�n�n����(�7	&��+����"?��{�Bj<$A��A�z��V9�����Y��U͵�� �/l��i�" �Ob�:��7�%#�	�/N��hV!��ھ͐OM �;�����,����ʚ�^��Č��]�Kr��~� ���B�f^-Q����;��c.]0v�Co2�]�l�S�]%9�I�n	ނ\�N9�%0�t
V��zǘ9,欋=�⎪jdo��N=��m��k�0�C?�թP��5�?n�X�g�ي��5�Bj�L8X���T�?�y���kF2%�ŭ´���e(L��S�l������:xI�s�G!�'�B˶o���|�%�1����C?�6{V��)+�U0z�)ԅw��l͖�[�y�J����4�\6�S X�5�@.a=��{O��w��m�M��	�WL���N`��h�����E�*��Z�y�y\.g�X�M������J�M�_Ӻ;��6�1΀j`��pj�uai��ς�pQ�xU���ӚNDR
��g��x�#��$q;��@��<��4�# r�L5^������y����b1 �9��W��%����~B\�G�X��=�䷎i�k����� "U�)��mt,�\�I���(U�~��\��S�b�H��5'�k�Rz�@��k�dTP#���S��y~�����l��sT"K�ң����Uϕ�X���7kH���p6r�^u�ASw�Y�@Z���'���^gg�#�kr��)���r��UP��Zu� ��ZtF35��7C��p-���Λ���#TS������"���c����b�3�p��o+Bx�=P<ծ�Nk�+�L T�<zFG��Ҳ�dq8��A� ����� ����)|~Ke�X��mco�f�򉃺�F�	�@��\S�ĵn5��/k}}nA;���y�?6��O���F2�"��G���P{�(��ݛi�B�L�����"mM]����h��H9O/�<ϵ��QдE�q�W�_wC�#��݄�|���@�`���'P���
���EO�,7,t��+4��
���\c��t��#��s�ȇ?{[7��A�8$��}�����6�����uA��8�}B6�_g���}���1%G4c��9#"�Em��`4��b��|�S,*�<w/�n�)��7V+Z�GCzI�����sn>H��C��<���Cn�|Z����?�h!gV��9����6�C��?Έ��O
OT�fvzB̴����b�@���y)�y�v�O�-,=��5N��t�L�|�|�e��3��'oN��ʪ4�bj���2�u*�\K�.���2��?��ٕ�_�����Zj�&�p��P�v�}�{�({�C	kh�$�B�1�Ts�1��~KNu�v*�-���d�nF���@��	k9�7]h3�nOr����LK{sx��
_Aa'��)���ZM鴽�^ۗ�jރH�-IQ�3a5�r";���(�D����kR�ƵY��6E�	�pC�^BnP�Q�ͽ)��ƹ0h��xڜ�w�Nl%��^�x�C�h2���V�}�:~/�./hZ��	V`|{�N+h����A#+$+K��& Y�g�ԮI��2�z��+��
IgJ�O,�c0�[��h@l�1�v�`u��(�(�g�2DO,+��N)��G<4ϒ�H&{���n��7&��U!G�W�벮�<�����*�Wo�ܓv�`\H2T�O���U���wk ���p\��&Wl��l8ی���W/��*쿀8�c`d��ٍx�4������u�s��$�wol����Ie��</��jh�_?�O��r����Mz;�4��lU�p�dO3y����m��/߫�%�Mgj^����\�kDJ��������M�C�AY��[����^E�g>���]xnJ��Ch����*��s��`�B���L�������Ǳ�W��`Նz�g�v�zV�����)�iI��B`uJ't�x���.n����%JK��]��$1�,9�q�{��k�<���z=,�ߦ�X��!���� `s��N�oj!��.dՂ�r���?�4Q��ȣ��~�K��HpQ�v���iƱp�Ќۃ���6�^ZGE��m�X{%���^'Y}*�,s��ѵ,~c��IQy8�s0gfvo�[��F��*�݂e�}��h=�
�HC]�	Q��Wl��w�Tk|�p�ĳũ|���)��R�E�	��h><$���4����c�~홀��v�W&��(��-�O��8�;�v_��,i%)�u��t�F�$8���n^nm�>H����+5�*�t!@��[A((�'5�
qL�7B��k��RE��n�zࠢ}��Na�%�@���BtSS0���t���ѓ��OO�f�����B�8�J����5����� iX-E�DN��z���q7��8-\��O�wk;�w�J1?iA%��/RL���?T���2d���T��ۏ�-�V�cn�����KHr����:�)���rA��t��n��q�U�����m�Jqa�\���AH1C��=#�<�K�(»ؿ�vz7i�o��*)�z��r��a���I�L�߾R&�����8x���0�l�>�&u��)!/�h�Ii�Z���p�B�[�U
ħ�~K��PGⰤDy� �[�� ��O��>E�s�,�'A�����0��,�0���{]�U��Ǆ�"�ȇ���h��nR��r�������T�Yo�~�V�jZ�f�s���5I�A��]����Õ����Om <�$���<���7������ё)��0�Cf��iy��-#͓Q0���*K��[VQ��޺cȌ�|Ӂ&P<���Ί0ub�S�$R�9�S��<�ՍL;ᆛRi�(�a��w�A�^B�S�F���Je&�5�dIx�x�>IM�F!���9:u3�9B	�b�W�Tu��sW��D��4�6�����\��t>5�;�o5�?����{���y�̋K�.�̣�~΅�A����W�6��h�\׉���d?�ֳ�_�$��X��Lh��yg�QU��.����!�\9x�[q�gO�1���|�A����v�*E[���H����f�(�8���F�L�ӣ�y;K�L/�kgYOMs=\T�_��+2�s�b�c:]�iM�N�UxO�����/�b�*xPH���a�{'��X�۳Ȕ!�00�/d��-M�6�O�������N3nKt)�=�uq���mIƪ�+���.�Q��s^��A8+�R?���r���������Y9�
�!#�m�X)���Q����[f�/���K풑Buo$�S��/w�C忠�m:�"x�?heT_uoYT�S��`�!����"�H���S�C�4�:)��b�C���!�� ׯ�du׏���R�)�q�Q�̈́�ʣ�f�%�o��oA��W� C��Y�vm�U���L�$�B�0����'����v!#�f�U�FS���2�P�E�9�|%׮[-؅��;�qy�}�C��ct6K�b2��$g5%^�|�8�V�.�p}eOO<�G ��X�K�G�oL�q��kE!�7�̥&䠹OB�`c��>���hܨt:]9�m��=d�yF�Z.�I����%jQ4��l�ivꔪ�L��I�s�o��P�-�PvLKd���G�4��L���7�壖��R?}k���d�~��w� +�����0�w��l�zu�H^'ih�'�G^��+Y��f������4�D�⨒�� �`N϶g)!�i��t�יqqz�|�j���IL�3H�wuӯGF�xPұ�91���]�)+�ZpEMfVvhb�gb��k�|P����r�� �Z  ~���Afui�Y�Fc[7Dt�:8�R�bjT��.�@
f�_����=����G�uE�X�NgJM�ý&͑{{յ��߷�YѴp�.���8���.�(�j��XH`n���)��W��^w�R�G�h�4ِ��/N�Gױ�Xr"���!\��.��j��Y>�o����IB���X�J���L6�����3n�
1��y5wOI�Q��S��4Mҗ&<ۢ���"�W}�l��h|#�66A%C]�L�sv/�P���<޲@	�@���G��>�F���%�@~4i �����ͮ'C��|���(G�0ha����}�q>�Hb�a=�=T1I���q:�ֲQ?b�ՀN������lE8�X��\lM'�����y�r����A1aF&<EZ��"z�{h���^e�@L��
�g6n�x����EL�?�w>7@���H�R² ���\t���9���C�͌��}�(f��ʭz��nd�~�7K�;��(��S�!�2������Y�a����*��]l�u`�n����AYJz��2q���LW�7����-Ne�+�c*��1M�C��_�q�x�$��%�즒yJ�Ijf�gt��>��"a�EPh������o�.�c�a'0�9]�|�w�Jۏ�΀�,�*������v�X�f��p��<t�:�Z�qA�!��w��<���d�0�nQt��9pV��Ϙ]���]���o+k�̳�?�M��`�&6$;!O]�ԑ+��-��ņ���������l��sO�&�iVw7�s���H0��zGH��B���V�b��2�ݳ����w0R�־�צ|o�i�|_nk�T����-�=��ۺ�Æ�#�%V�r�ڛ.|�{�2a7���^�&����@%d��k�e�/��@���f�<4����ᕡ��>�"��H��$š�]&�[l��-�\^�����R�eQ5��<�ʊ������:9�������R���V�� �D�6�d��ѽk�I��<$�҇�n\N���H��Scy��Ͼ.0졝$�g���<��"b����5r��q�<��f���u��P���Ķh�۩��:˞�Fb@gnᜇk��}�2z�|\�rf���M��Q,-���ى��˙:���<��K������/�,ɕ4��ǵ�q��Z1��G�t��Pm�s��N�\��Ŵ � ����3o�%�~}����Hj,t�)�*��Z���$�C�`���{�\q�H\���:�;��M"�k;������6D�)7��.��N����nz��ZPgM����9�Y�~
��ZGG�{��M{��������Ŧ�{bδ�`6{���[�F{����}��m��]K�����7VjZo��2�J2:Ԛ7�L:� ܙ�!]��\u����9^��#�����\*]mp�-X�������5騬8�3q����+uY�X����9�E�ȶ`��f4c]�JF��y %j�H�H~�&e�7j١R����f���r1#M��*�v��E���zB�9Z=OV O�u��Ns��X�(�6$@AI1��:�e'������3����CsВ�ǆ�Ѐv��n�i��7�
�ZJIh&ӈף��]t�����=ӦŠ�(�F�\eI;��,��C�%��>���!��� j��qtd��m����l�g+�d%�ߩ�~��}y��<DdJG�ɣVݾ��ϫ��l?�N������V�N]�-�Nҟ�hw!?C
��-��"��zO��0��8m�1�Bh��`��[-����g'��a&�y���M�����MYc�u��sh����\�t|�ʕ#X{j�H��m�Y|͆MF��d��R��\��蜸t�5g$�E����zƔb��v�5��'�a����n���k<����5��&�!�bM�"�1�s��	�_�沰�"���7��"�w�r͢٬^錗��؈z��7�wh��y��������W� ���P%�� r�*_j�-�4��)y��r��-7��PG��t
=>f�P맬5 ��渻�@�#@�ׯ���uI��4��m� 
4I(��n*]�78?Mv���Ły���ճa^'��S��B�u�����R�Y��]�{Hf��<#��ť�L����	�Y1�
�������%��$�� ���`o�Xx.W��&��.��=�-��p�m������"*D�<�`����)�w�<1>��C��50� �;��B����2�DˡF����(Q�3@;�Ĉϱ� a����Z&e�Y7��I6���;d���܅O�����[�H��va�lH����֒�G������������9����X���p4x3��j�Wo��>��
�t�*�Q�h��$�]�����s�&(��M��s�F��3�D9��L�1�٪���j��N_DoYUt���?�DR����7��~�Zts��e/E,�Fp-����f�@�Ȫ|���^�����n��WW�&՞,�d%�:�Q���0E�f{��@�pz{}��Ų� )���s��\RP<�W\�g=�.m�r���T��@�u>K�N�yW孭*bn��m���N��Z�T����C�$#Ǐ�����h�W��?W�n< �#�(�n+2��W�-P����D��]kR&N���Zh� �e@��}��Bީ��wX@���,>pƭd3�����4@/��������.�X�i����>�4�|w^U8㯴�X��8�@����W����ktOXv@�4�l���"1Yő�>��{������[��p��!�Ƙ�Á���u3pߍ���6f���S�7*��~j���T�u-���M��#�(W�4�R����J?��@2��5���������Ԃi��	Əv�\B#!�	�T�SD���+��{Kp ]ڽ	{�3�CY���:L���u�E���_�������H3>}��s<��*X�)˕��\�:V������_����nwx��t�Y!���\ҐMz��}9c\�U��y�ǫ��~�#��ч�ﺕ��s��2�1u�FFΧ���lO�����D�&�ʫU�>�@y<^��i�rL���Ȩ��S>���4���!
�3���%��^c��i�k��!B��L<)"��r���YF��6���#C-��[��F�k�d�i�_c�[�c����G���}՛3p���πg{���d{��	�����S<��CVI<��!��I��o�Q��g�Rni!��7�E�E�`�,A��cA1��,�����9]��*�A)�t�smV	pr�!V��1}�����Փ*��0^D�g�q�.�N�|TwDF��*MT#o-{^��h[���˽�Z(���
�|{X5*�E�_	I���+��&4���-2�6}�*/K��Qu� V�&7{�pY�#ņR��	;����o��k�o�Z,�[� ��Cfŵ���/��Z.�B��I��̛r�6�i�?
#��j�?��>�([�n��=�q���10ۓN�o�x
V���P�-n�|�np 1E*�%Z�w��t#~Ki�V�E�R ����_ɋUW�����j�h��0�����t�ztL�yy駵���qL��'Pe��sԜ��Q~��r�{$���W�9�ǯ���5��R��ŗla/%U�變~�
o��X�V�-�U�L�k�{��?a�K�-���r��Z�L����RU��A�9,��1Bna�?��O�i���c�͞I������6�Mel7�o`%��Q��4����$U��nLRz���2���G��i�w�̮Չ��8��P��^g�#��������w��I��ʔ�~�%�BX�{%c���X�+·O������Z�R5���w���4��8��?��ُi�%���Vd(��~=�MS����&�֮�� J�Yw�Yx��kt��KA-b�"�',�e��8��0Z�	��H$�РLQߨ<	�dh�d4�n�w+,j���Չ�QL�����������Őy{��l�an���jJ)W�7�A_��-�T��(�	�Ļj��a\� �fS�r	V9z��%��#���p
� �R\��G�v�;�Gm���o���� ��������I.g�@!3/N^��0,�?�O-�����͡��.>]����C��KT���Z?��j�>��ݻ�C�� Ҋ1��5ڇ1��g �"�O�@ qFYe%�Aam�^�P~ˤ۫���|O�v�%�����y�o�7pc<j^�F}�$�|��\ս����}(���r}4�Ѫc��q�ƹ��!��c!Z0���Q7*��.����0��#�-�[V�#�j��a�
�MJ�GY���x�/�,�8Zk��d6��j��!:BuL
����p���y��]2>���kA�l���<<��.����+"\<�{��b3�P��?<����('�]uW#G�n�mOf���]bE��w������Å�|�wS���:sĦ-c��XD�ү�Np)^D˺�ؐ:����i��,����V��tu�M*��?���o�-���_'�`�_˸ɼ�K#>�Dhv,|��.�je������b&�W�}9!!h �$f��h��l�?�|�g���Ag9J֑ϱ��wFq�;]	_����3xMk����`>)�#���<��ʙ"���1	p�2g�l#0�������d���(Y��eCkn1�OQH�D�Ó��}�@�� 0H^rT�O���V�a� _�Gjβ�V�4��&<�I�fm�=���5��}}���Z��@���>*��k��uJYD.1��}�mN�\��*�aF�K��.'l�OyL8;{�I��h��xhv6k���?��֍��$#Ȯ@TGbB��-GTyp���ݑ�!)U��c����O@M���B#W�$��Y��@rCz_D������FK��"�U�g6��ܱ3mr�-������m�|$S�0��5�Ji�]���ؖr.F�b�y>�}�"|����*�ޒ6e�?_�U| ,����z�X�}ܟ]� 6޷(��g�.���̇�����\�+v��x��:F��6�)��;{2�]��l���Gy%g~{��gC!/30}�e�_��-;�S���|���V���,
�-TKg�ď�B�����C&~�љ�K�Φv����A1�,��`����k��1�o�(A�0�	`�t喙�"&6���7��󑗟1��
���1�Ɉ��;�hVK'�Z�GM? cnk5'Jޝ]���k�Sȹ�3�{!�����d<�~��X�}I��o��A �а�r�<Ш�f����Z�8��A6�Ѱ(��c'{�:����/�Փe
�^�����yKo����A[.!����4��8 �k2&oN�ST�J�gU��H��ױT��Fe�=���q�*|(@`	�2��[o	��t����	�Qb���Z��,V�*�V`��;�d\R�{gm��u�r��8�q�/��(OuH�n��Ơ�A�VԴ�uJ��/s��*"`�B���1��)��e���{��%�$Ë�?��oBwŤ�_��N`�l��Q���	6�|Ϸ��5����A��8S��K�I �֡�Z�1y	�w�}�G�f7��=��� @���|Ny���a�4R�U�1�����8��n�ɪ}-2�!��S# Γ�P�y���rL�J��{W\{ϪS��x���U�n��]�'��s��u4*B�E�\c�.1�����؃������4�ҍKVB��x;�C��t�U�H>S9e�Ԣ����`kfsk�n?��Y��My�v���V�E��G���a,��{�i���9����S��q��}ʸ�s�ܚ���Ё±�@��tf?f�_���mZ��hx)g��v����p:<�&vqZ�ˈ�����1�H۵���T �sڹk?��5��ע���Q�wx���gcC��1̿������-o����O����ʽ=8�+=�k��"s�=oo�Y��p�=i$��l�	@]}���v����(�pŸ���b��h,ҕ֩WSD8�>v�Uy��7��Ax�20B��+/��Sr��|�b�TxZ���vJ�|���+��z
�������z׼]��;�/��%{�4tG����о�l�u��H�!�Uz���U���J�B����TlOE���<��ToI�7>=�  LT�K�I���Yl�?�M���r.DWwM�b�Z��<k��>[O_{��B��k��zR��NP���g���><��f� :ƫ�A���Fb(��{R0��uۚ�p�Ǖ�f��c���Y��վ�C��'�0
�`F��۵�/[)�-i��yo΄���k��G�����$�D���EqD���S2����R'/c��ųT�����T9�^LsVn5���,+7��J9䦽��ty������4 �
��ͫ��h����<r�ҥ��y(�f��7����{]��f���B��7�ȡ-��p��Ȥ�ʟ! ^*�x������V*�*A=B��*a��Jʫ
�[��!.9�5����Lܕ�a��70�q��d��̾g����+��l���5��fU��r���p*�CF5I�`�����óH+�ؠ�~Kl#)�V���W�Mx]��*ϟSV+T��a�a�c��
� ���W����o�a =����įz�����yCz�>`��y���pړ�H��������5�O"��Ւڋ���s���T��^�I!��ў�vQYi�i�β�������u%Ex�:g�����T����5C�S�>�T-GHOP4k"l׬��pu3��)��7e&P��Vq��0�>���@ޤ������Θ���[>�Y������H�(�T�N���GC��l?_^Xa��:���6��Z��{��s ԋ>
j��l:�2�� �>[n��"��(�����#���-&.�%�=fz��^��w_�',�ls���4fx�:U��j�(�SC)������(�(X���(�.��<S�?<�}�U�W��HuU�$��m`.6~Eҝ����_;`5}��%�)�_���/�#����cp�FY���Q����,��roX�T��_�	�%&�p����J.�s�F���r��ڎu���X!|���S�
׮6�K�g�p�x����Nhh���;���?�M��Ӫ;�[8�Tq�h�3�-��5���L�gMs?L�I�����Z���.��ypz��zd7fؗ���@�,/� �H�y��m��Wd Na@gj�
N�5��E'���'�a��+,���>�P��_����}�D��~�/��J���AG-v9���7���m-�f�	���B8?ߺ��<������9�t��+|�&�G�2P���"WI�,�BB5�~��>����sFGBm^���?��t~�T���Z���r?|���.�{����6
��<�>=����^�0B�KL���c|�G���׎��jL���$H��ie}�T��Qub0��*Fi߉Y~⇅��"�o{�f܌ϗ��c�o� x|��3z4|���f ���N�?��b�خv ����4��~	��Zט�(�������s�^����K�1�^ t����D�4Mh	p�����k�Ӿ���^A�Ty����2�JSn*e��ʱ5B��}��� 9���X���켛������������4vC�����%��NF˴vvY��ps��
[��*�`c�PCr�k��r�]x����q�!K�̴��RHb�>ՠ�4�(i^h��{�Sn^�_OB��N]��|�dZ��2��ēC��ՠ�!H��;��v6����i�~W��Jׁ.`�A&�'@8;�g���I�PLX9���%�&o{t�8X!u���#U緲E�I��`�f�N����1�'x�����Zmp�0 {	hxSF2��;a����s��� Z��j�X�}��#0{���15��_  ��RD^J�U�]aj|�]��
����z����
���=�,x����#&�$��zc�p�kZ$�+v��&F���pZ�0[�Ņ�Vэ�樯k ���SQ��(fD�#��/���n�ʥ]T Q�nSՔ-��T�=^��TQ��l�^ʀ7�8l��V���XX��P��@�Q�-[�e��= �ݱ���J����'_�)�z��.t����Fm��Jr�� ���S�\�c�00�%�y݄�JHI�et��lQZ�f�(���k�j����P�Mb3��]�J���|R5�<.߉�;�Ta?���Wގ�;�*T���^O)҈�p���V�,V�Ҹ#�hXiG:�/FW@2�)Į*�a��[���3����nrq�&(wG�Y7�C��O>����;�
�I���kXdF__<�9dn����U4G[#	k4Фc��ox����'9���mA*+�¼�I���y����N�:�6�;XJM�4�59��|m���	#�S�gb�'F3�S�.���y��b"�s�*���o��/��<�i���R2`� ��8_���C��gc�#�A�ܓUj`����z�FB�3���{!��݊�W.�>���?�1-�<?�8j��0��$"��IL�X�%T2�l1�,�����]���P �s?<c�4E#���e)M���m��q�=����1��	q�-8�_��n��n��7|0�C>���d�nr��q�;�:� *��?
��R��{X_+Z���'�.u�=�tӳ��q(f	��?>��t`^pX���5�U�c�H�� 攰��7��̮~�WC��mx�����z��k�aGt�,�K�w�!1�,<{MkD �l����x,���=��Ɛ]I�4_�����&औ�z�s3���F���+�s��7�u���E�Q?DB�Jh\Á����w�5���x�d+�F؂��?�ʋ��k�����>9B}��'�:��n�_�f�L0׺L*3?O�9��L�̼�zi$�B%�(��٠b��s���j��|��@ٶU.�K�'?�d|�q,�\Er��F�Z�p���
h/���8�͇`A4�biv&��},,�Q^��Ϊ�*�9b�Zș��?#�͐�9���X�B8�[}�{sݢ�5u�Os���d�����wr�L0tC�z��m��JAO�_��d�D޸��l����@[��dQY|�h�\��P�]B���PB�>
&�t!h3R��_�j.�d|�%ثW�����~���!i_+�C X�ط�A�j4�#� �t}�b�bF5�r-S��j�����V��D�P�蚭�X _f(��%3xQ^�VW⭅����VG��÷$�0�h�ќ�������;�#V/hN�d?/�T���&�E�Ԭ=����r7��q�H6�g���������B�dW�R+:��>;��t5�?�I�̽ς������p�Ug�]��߀�N����NO�bѵt/.}?�Y�!�0]^ʘ@��xI<�06J�R�=���#b���2���JX�)��%O�X�:B.���O7�s\�oz�q��ك�%Z�=jj�-BUe���i���\b��_�?e6k���mӛǙ�=hĲ%Q�/�-YY=&Dz�� z(��)ҳP]�j�"�����/��{�T�k���#n�U��8��z���vѶ�.�S3��6�����1�H�bb��`� ��h��i񇡶6������Nu��#}?RDNչdmX]�{X���m(�<㨝����ƽэtxpH���q�Lb��xB�E�_r�^��/��?O��8��s���"y4�<�"+�H�����X���3�����va�~�>����Oh���>�3������͒�CzT�I���$?ZeCb��εEZv�=)���@���7UZ'���ƹ���V�w��u;�lC���;��A��`��̋�f�
�� 5�vP쌥��2W�*->��6�X1l
3�]�S�]��B���R9I��2">��>����	Ef �4�K�t#4
�[��7uC�)�n8ho�U�V���	���m�舨 ����ҥV�T�[���e�O���Ҳn�~^�Q���	t=]�V�5����;f���ǩ�x��I�l<P1@T�[� ��H�]C����jI_a�9�����\',Ry�2Ō��|R�B�zf4,�����ӯ��W��n�y�o`*�P Q���	1�!�n6@具XPR�F/`J6�� ���ꏩ2nT}f�&^UU��;��lpĵ��Hr]3Vg��o;}��9:ӌ��ؔBQf@�ib��@��Oc%!>�s�}���G*V}����]؎���)>:u]͇讈�^�h$ᅝ��� ��t���˙�\{)�;h��2w�({���+7��Cdc��?�o���c�š�N�J�����b�Ԙ��-\�'��T?�d!ZUI|�����z0��p�zW�k9
`в����ab�מ�^T�K=G�b����솅J�.���h���"M�Ȝh`�1�p�j�y�c�������\f]��@�6]cq�j���k"S�\e��#��?�$�����Ϊ�b��Բ��*�B��2]�/"ڒe��oLi�*�7�0�5�X�J��s���WE����k<�l��q�M#�5��}*�d����LH����}�	|�������@����F���ugx�}�q���A{������&�)z{�c )�a�a/:�VX�n�x���ZX29��~M	�`��L�ք	�d�
 Y�J�'�^+��;���dL�-v�:���ԉ��8��w����
;�GJ�tC���Z�Jec��x�Ӱ��n$��i��ib_���b�����fc�E@�E+n���:����*�|]�^<f[~��A(�.&tĚ�A�s�k$��[i�c�q����V�7$@IPf<��z&�L]��x�w7��?{֨���gr�Gx8?���u��&1ep�c|5��쑑^2�*��uЅ��h=Q�1�wI��X�֔)4��#�I�K mg�J ���D�к��E��aA;^]���F�@�֋C̤��H��d0���U9A�Ι�D�)!��f��c���a
���(I�����Z�u�N�g۩!$������n������ࢤ���� �E2��Nՙ�Ӥ�	6K5�\!�a�W���}X�x����sw���X��Gq�#`����O�ֈ�0_@�*��aI�ϽP��sSB=���3ģ��)�2�6l��y�(�-���"m�*Iy���Z���D��J�O'��%��i�Z5G��D]�3�>h9M��O���U�u���N+d���86���^z��ʮ�ͺc�$��c���A���w�=e�b-k����E� ��}(̨�vt������`kYC��s��?17uJ������'����`	�_2�,����'r|��׈�J�N�i�匥�h�6����DRUXS���<4������y�!��{��N�@O'�f�����ґ{�ԭ@��3��s�D��9�8��m���.��GUwk�����VB����J$�B�$ƣS0��x�Rl �ᄕO�f�����b�Ct��H��./���	e��lmcbwO�N�n`C�	���i��;�BYS�'c�:b�}#ę��n��B�ܞb[�ID�p"��	�e��0X��aZ�,�dJ0��64���\�ҧ}Q� l�a\ڢ(�Z�Nf~�<���*�-�����n&ᣈ���a+D�!��$7��ͭF�_�^)XIRt��Ϋ��oQ�w�T�3�����"w�L�
v�t:�Hi2�C�r�eT|��-CB7B��DKD9��b��{�B��/������H.S:����uݤ�z/6a-M�	�|��J�M_7tF'���.ψ�4+�,���VCm����s~�m��@�Q%�T�beȳ��9���Z�n�(ޥ.��M��S��b�jD��|�6��nx��a�N�"��!W�|��'b�w�zO��h�)��� 8un�����Q�}㗊��F��	��CE��h�����s>�딐O��2s*��ߛ��!��<Z�C�� 7F�dL_A^��K���
�Rd���K��a��<����
�jr�Q��	��̆�f|���W.��WX���=n�˙��,��ι�D�@�3l� +��L�s��1�FGᛒ�y��_P�ʗC@�(w��]������)�0E��|�_�{�#\�_P$=��hk�����oÁ�_�,'��O����-K̼�B��&g��h;A�&]�����������~ ��Dha3����<�KK�RL8k����zk��[�����*w)�y��>k���C�$%r��9�"��^� w�%�jv	�bԭ9���Ŝ����'y}e%_8�l+3��J�͛5�� ���`��l�)�:�z|(7���ɴ��\lp/쩃O����ג�W���U+����D�	6��')�EZ����U�)��V�AW@���w�I^d]m�5Y�hPQ�V��s�mʬ�/��#�-i��R�����Nu���b�j� �gV��u��D��c�y�F�D�R�E�����K��i��Z�Xh��$tD�����$���?&�$t��l���iD)1i4Қ;�WS�oU;�������}�MCL��wN�I.?1����,b���Um+HЅ���Y����.�Yć4#����7ua��.��]y�?s"��6���|vx�h��|�T>�;*��w�C��?�'�'ei���e4��	�_��b��D�,c�sZ���sȍЩ��`�kb4�Kr�U�bo���׭�P��4��r��e��JG�H�k{��ޭ2�'��F7���n��- �-`��
��	�O�5�H�.�x܈'��*��^sq�~Ĥ�ĿØE	�=&�^�F� ϹOܹ9-����:�Jx=e0l�@�*\�m$���mJ��	8İ��
³�(C��)t���t�J���Z .�H�w�"���b��Oc�:.gKj\�9:P
�������/.E8u_�Ԡo���˗�$3&~{b���*��?�'o�6DWRKGtM�0�BgY�:N�2��{X�9\��� |����|�S�r�.�9oZȟ��s�[N���MDȐ��5�`ȍ�tKMp�M$:�>�$2�����ӎ�dh�`���4��+W-��Ӿ��]������X_��ϙ�T�>o�[���r���><o�\��jɍc Ls��i��h<���\��"�K�Y�ܪ����r1���D}l�2�����L���������E�T�]?b�8�m����7�Z���\��UFtL�x�]
/8��X���ȫ[�F�Z������~�z�똀��9H��������I gEYWJ(AsG� 1�t��Ȣ�����!�KkBN��rlC�C���<~����@o�ᛢm���|S�V��h���w�"�_��OKQ��_�T���L����Z�J�4}@�{\��{.��p}I���Y��e~Qc�ѣxS��{ |r`NO�D����4�돢=����źq�{ex��A��u�1��?�ϸ���.>L[���v�+���`�u#�=���j�I���I�w��+��pK����0��%VZޥ�TT���{���42�kt 4��V�2���C�_]K�� N��P0�9 f����L��y�<�=�&��q��x�"���_p[�V�U��ַ�>qXG|wu#�J���@"8��8�$8۠�T7�g�f�C�d���qޱ���(׈r�Q=�g~N�F�W��c��Ul8g6��Z��L���f�!?�ڽ��u�1��_Ѷ�5��yu ͑t	s�X�MU��ڊ��j�u+��/������R��&� Mu���ySH��M|}��f_-��%3�ϛ���'~bRȬ��3z~�.��?>�M}?`s�.	M#����- $��ӯ�$bM�x [�ӯ�.��i�N�7H�7y���[9}�G|�N?Q��h�^��tXmȰ�-4�c<�	˞�~�8�;覨8�o�_j:��r�Ԍ#��������pY6]HV�jc�&�$��Ӛ������l�L|�(�ֈ�3x�T�r�g]��R�t�����E��n�֙��C0i��i7:��N�d=x
�k��׆<�'�|QQ?ͥ�.h��;�+�P��)4��﬎�p"'�����Z۳�����^�炀��kG�X����,�8�
;C`�;X��Nc�Su�K���.�՞���5�J P�Y	���5t;hN�X-�fa!�!���/K�]@�OS'?�+0f�:��L�ڣ��0�yA�E���*4�+����,,Re�9[ǿb�>	h���k3mѳ��ʵ�WXށ�i��WOG�$��g!C]�*���ޔx^Z���sw��:��9I�5������������)R\�/L�Ά��9���H~e|Io�d�9�
�_Q#F~��y��͖�G�UO�N>�0� D�ye~���1�A�pmL\��xeLr���`�4]���Y��s��dsZ��?d�����oa){� 
畀��/�=��C~�6�}ȱ�"����x�E3�'��Uf�>����"�D�k��ߞF4����{���'����#]��3�^c�|h�8�ڠ�q����J� �!~�B��TUjkQ�/�ol��9׀& Z����,w<WN}�
�''P9���/8�d1V*&a�O����:_���9�hCQ�UZ��i-esA�ۊ����&ؒ�3�!85+���yo4�kZS��"@5�hǶe�V_�
	h��w��q�-A:�n�����Q&z����T?鈭������VmUg�!7�+ݍ���Č	:��j {g�x�.M����k�޺�zO#��?!�{Q�Xчc�42y��Sq7;����Fu�~O��=���=!�G���*�6���.�tx�����߄��?�r�H��x��Zc�R���t�:n��72	�?n*Á��Ŋ%���Na������߯
���'z�/fX5�D�gM%J�M�g��|��l��s g�p�bP�H��?��.e�h�����
 ��ίe��X#��l�LF|�e%��ל�fH�j@^;�&���$�
9������+>�8@8�f�vK���3�G���ʈ�Ԯ�f���>}3��3)4,%��p qCb3v��C� ��ۣ�ƅ$������g�����c��E[Ey�0:���T�}·/���A4!�f	�_�)-�#��޺�\G�x/��S���P���U�[�ڎCS�
�s|�
�-�{H���9hE��H�����z�e(Ӵ�F{-�������H�35.-XN��Y��lp�h� �G:(��lR�����E�S
7T(��J��I�m��A�}�в�8����cr�ا.So��eR3>��
�4�
�_��2B�4[!"�権ɓb��̲\J�+�h*�s7 ��tͯ�/Ӂi�j�# j�H*��A>�\e�/����E#��itm���n��/\��|�b��bE8�k�k��>vz�(<���pP�9L�w���,\�c(R7�)���t34��vn�jxz�2��y�Ms����6���3��0	�9�m���Wt)5y9[�T �b�P (��DS�����]�9�0< �9�-�5���2�L܊�ؗ��+d��ܿ"b����,L�ӊ�4R	���B�	u�����bC����w���Gⱓ	%˴�J���ȶ� �̡��"\( ��F���͆��i�㒲��A$֟����s��l|!wX�Sy�1����R��#҉�i`5r���ď����	*ԣ��hkExd����C�kt?˰{��C��P��	�� ~�H�����F����FZ=ˣR \LyF�A;q�O�TmƯ��TiMGl�yXM
�$2*�AzļGʻh	���I�+�1�[_,�})��""����_���Ӕոo����{>9�+�+_ڪ��B"�1�1��h@f^���s�s��Su���k���o�>zL �o���l��m�؉3��پ�ӹ~-��܈��Y��m4<��H��3�C���}K��¦E,5�t8�͗�����l���Cl�r�#�hŏ~��4}^7a��Ý��I3������H8�O�\2���Y�Tf�t�t/¤(*��~��J�Y�7 !\���u�4�8s�T�ٌ=j(����a�'H&Ff���ꌡ-�Vf�z��o'0o�7�#.�q�h@���9]N��*x�8d��\L
�Z�bnS�j��7�p���Cq&d?LX0�9�g���t��cR{��G�{W:���]��a��,b���("v�<���=
���O�#u��wY�y�`��'�Z��+�c��6w�v����q�ި�`�\������
u������)�肵����W����w���L*��{X���U����D�=�or����������	,"d5�ROP>�R���7�c�{����T�۩&�tt��{k�Sj���,��xz8�W
Q�*��\��+����[����Lb�1|R�?�nB'!��o�Y���r�*0�o %��
f�ж�7WS�p�ZD& ~OϟU�t�*:"�K���Wy
�K[�J0��F'(Y5}-1zH���G����N��B^`Txw����g����A��I+��_ï��֖�9Dy-E�?��ǫ��H��1ҁd^�Fȑu��b�������G�S64��4�c�K�^~����q��mz�,.~��r|)~�p� �֟�����hzV_fbYƏ��WzbooS�ʌu���|��<�ջ�Gp~�^�䞶���:�˵�76�Lb_�-�<,��^֪�x@cJ�*<�@@cT�O`��n���;):
���7f�]&�>x���ƍ;_����B��U��9|��y��E� g��g���W��Q�v|���Ë��XQt�*��Po�c)�q�y4���oB����el��pJ~��MK�K4��4���Ѫ��XB�V� �����Z
K�E���-΅���i���^��@�����`%���$qS�:����M��Y�؉��R��.R&>Ea�b/<����TRn���,�.�����Ỉ�!�	��2Rs-h���6{O���o���ܝ2ǂ����y��V���1&s��e�Jϥ���o�BʞH�������(T_�s�@z��G)@���ͼZ����u@�&�"m�H�_>qx�wS|�ر�="�K����kN�c7.K�3eU�������2fۅ��6������VhP�T���Y�r�G�P�ZA���y_C�I-,;�˲'�3E_���0�ӢoI/�mS���F�6"��	�TK����$�_�����{�:������*~�J�K�\"�v'������Sɔ ˵�����V��[!�7����闏p\�x�'W��vG�6EH�4QW�p#?��s�Db���
�T�q'0�
�Ei����B�PEjڍ�����q�s�qRJ]ψ_����n��Gf;�	��r�\�CsС�ܷN����0Ûa5}֓����GNM��r��*���Ă��oȾA�w�V�禆�Ʈ��r�J��[꒟���>����!e(����W=��̸~٣8�/�����dJ�ST����in��=*�S�?#-3���qj'�9��>�s�7����A�Z�������}�3ҢV '�X*a(�_�t�LqʝW�2�!Z��#�K��fFy�J�U �=?VG+��|�%9�����4P���*���"*T�Q�^�V�*T������L���i��=��U�=�s����.�:� �����D9v��g����+"�Ӡ��;��Y�rZĲ��t!q�
PBSƜy�2,�=�n����~���o�r�[7X;�G�"�P������h�~�}����]1A�\&vt!(]�[�cCB�\�]�	��� iɯ.b���|��h޸ �������i3u�	X��r/��jW�O�p �H����N3����/�pj����˙y��j]tՌBaa����i8X�	;j~�
�c�Q�3�C���ٴ��n������w��<I�-ے[%��=aX�|��T��R� ����m�]�y랷�y�2Jl�Q��l����4�����
�ʅt�P�j�*�~�l|6�)4�N!�U��rx���j����̄������@�ꜧ��e���=����P5`���	7��v���G~p�G&��x�n�`�;���i�������_K�I�q}�ا!~	���]�\�=[%R���_\{��%B���!B��ID(��#g��g�O�O�2�"� linRD�	V�p[5p��M�}5H��8E�-?Y���h-��W�|������n�X��}�A�i'��j�����d{���3�a�A�X�~rj��F��QT����2�W�w��7�XX�2$�\��/�[m^��"��y*x���Os��#����H=�N!���a���w�D7�<j.�xi9 A���&�\�4��g @��8�d(����T�T�i�.8�_qO�����tk�S-�d�d`瘔Uo�M���I�����7.��m�Vm�L;bX��o,A���K���k;�F���b�մ���;N���%ߔ��eR�}��@�YͿ����D�ٛ��;�F��lQ0ָA�!���@�V�%���tۣ]���C=�1.L؞c6hdᩅ:�0�ˇE�*�&r<��-��=䭗�.��4͓%��_g�շ�eI�����]^� YXUA���n���l�b$}iՂh4\���U�)�X�uVh},R���<h �#��A%_T�U7��\�4h(#�2�~<^ {�0F䉵��Γ�Nh3f��k�p��`��U��ў#�إ�:KP\VD��u)��:���-Ju&@�6@$�r�X�r+.9q�g��¸U�sR�e����i���om���}��/j�W��Ԑϯ��G�mu�i4�8*�V���f�����e����DE�Pl�)�jЏN��.�`C�ְ�ay���/½T�qZ�
�zL���2G ���Z������t�p~
� G���e��o�q]���6���a�6*���s�� ��������2Fj��ʗ^�pn}L�p����a��ذu�����c�@�3%��d7��:4Y�u���d0M��v�����d'o�2���^u��s��6� �[�&[&�hҒ�K�.M�K���a�B&�����v3���y��$~k�d��	?�!�_�
n�״����]A�5�<�痝���+z@�F7�?$5k�wm�_��^�&BH� �OMF���}�Cnb)�"=o0l�=ͩԾ-)}d��"طR��d�>O��Лo���E����	�#?�ź7'�/2	H�:O���Wz�sId^ �(J�t�C�񩙸���M�]�s�����˦��J�hFKo��Q������'�w��0����r��c��Z����+�½/駅��������(���W_]ךs1@���`R�1>>�=����.�����l�_E�q��4�~ſ��q�������l��m	���.�cJ!&�!�������m��C؊��[�f ����J��kXGGҶ�Is",`�W&��Q���.ȏ@.���cԖ����|�����g��y�IQf�ĸfCV|�n
��}@�D7:��_�/&N��`ZP�z,9t����K��)�ͺw��MW�66�ͪ�tݾSH<���x����쉍�f_�{+T�x��%b_쬻�_壉lmղ6Tl/��$>I�NZ'fz�S�
�9�@�g6Db$�\�WُteccF�Q]��3v60o��b厭7M4��7� �>���%2����u�������_n�es���H��,��}@�#���Z6��l�%d2Ά���Hk$3�S�<�,�VBJ�^S�Lt��."�/Pp����J5��캓p����hѣϜc��hԣ{1�L�L{���?�㠁 �yt�3��טy��U���U��ΐ��ɰ����N�v�Zr��`)oE�y��E����$,��H���|�4�5-�g'�s��sd.5�1�u�n�a<�����g� _�h
y�jO]MJr�\���3��,���Fy	���h^��	"��e�������K7e�3D���ĭ������eMz|>����z6r�~�u89a{5T�!Y,P�Tz6�e��o�])�e�&d�p1�R�dG�A��!��M������r�KE�~�e���ѣ����h�Զ�^��Q��):2�v�'��С�ݶe�x�_�pa�Zsj�a�:.p)�q��E�/;c�i{k��P����1�A�s@c��0�Z�!����A;�-�H�4=ordi-�������jl,i�dt�|�WAg���MSkZ��Y`*%,�`����R�����.1�T�sl|~L�=�9r"���z\1B�C�Y��z}!���[���iI6�_7�7q��jqLDm�1v㶗ޱ�MTu��z�L[�� ���h���J9_� ����<t;���TB^�w�
��M�`�S|KSyP\�{���߿�iMd�^1��_�b+��\1D�1T�Z�N	����g�==�d�sC�v-՜��̻}'_��y�B�Ӡ��ֿI��j��x��J��'�e�ˮ��ȨL@�3T��o����)Q��J��x�mf��Q2çT�.|��08����_ ��&F��L+1� ��77dn?���ށZ_��8|H���NN�d� ���n��]׈A-����=�k�
p�Z��R�̕��|?��F�1?�e1�� �:�v�12h�ù������x�?�ON��UA-<�U�����d�Dlg�]3�m���7�xz6��kb���fglQ��cЕ��D��<����&L�.ѿ�ΊҨ�,� ]�<��D4/�]p�Ht������b ���gp��Nӎ�4�0�� u}Ts�����̏�b�X����ܝ�`��'�V}>d(���&�?XV�+�^��Vb<ƻI���	mOeAm��+�.I�\���;�'÷��� .z>��U�<����C���K�8�V�	�Vw�:�$�1Kl=�ռ�y�;�2�Z�_Ylӛ!K�#ܻg�����=Ϭu���S�aVo�fI��꺫���좆z4=~^xj���ƅ#��[��A�荲�)���!�5��Ŷ���sX�%C���r��K��������V\����'c�U����ʣv�'{xtd2OY�&./U>��i�[��F��(%��/z,��Dw����Ӎ>�d����:�TT��83o�kǙ�����Jhj��a�Sg�W�Bh�b#��� �y�2ſ6%7*���;2u����C��O�d�:lΗ<�cW�[�k���٬y۰���{�"�@�&*����|H���ScORi�3�6�v�Ȃ�^���^�G���:^?҉�~)���܄Ϋ4����"�$�7�=<�h=)p˿����
r�⥘�����H`vmW<��N�7�i8>5�&6ĳ_�	'��-OE��fq���$uY�Sd���Q��鋓�.�����}��O�:!�n�a[c.�ܟ�~���n�Oњ�͞��w��
ѡU���gRZ����N��j�v(*Q|�ƞvv��H;w�,A=Ɂ�~�[&�����Έ�)�6ֽ�V�4�(�˃��n@&�
��n0G>��X�y7���秶+�pUf����(�X���;\�1��#�޴VЁ���[�-�b��*�<f��gA'�
k���E��WɑI+3f��pS�':�;�7�����K�8�~�ǁF}��P\�iX�s�<1-]`��p��X5��幄%����g^6�#���E�FW5�kx?��"�[��R�/ ��Lo�-u�{�}�b�9����#��~_��2��h���c���C�U%�=yŪvGb�ɫh� ��c'�L�a�Zċ?$%U�ñp�3�)Ѥx��m�����HUSx;.֟M�H墕�h�x)ʹˢ�=c��;��`��_������5Q��%<#�B���w��Ědz�w].���[�|�t���Da϶sqx ����Qܧh�CGM�:[	��B�,x8�
`0�ͼ�o��f5`}�j�&H~���8r����>�mOa���H�8n�����"� �89V'�!�?f�E(�T*�
J?�T�o�B��Ш�h0�����0Nxf�,d�)5����{�
�G%�q��?Y��a���ޯ�vtVPH�єUZ��O��Lҽ5ל3�iQD��s�Ճ���ZL׃�Y�A� Xޙ%0H��:�9ת��D�����d(��8���O�wY{ t�`i}�Ë?�b!�F{:�0˂D�5�)AVHx�k��o��hhT���*һ�୎ ,�K8�y�-EX�o��Ю�J%c��#��O�f�y�O��:�{6�_q8m��BJ�1��D��s�=����R�/q��6^��ڒ@���(�m�[�R<��7�9O6Ǫ�FR`6�jk��?�Φ֙b�%w���GQl�aJU˔*g�1�*H�^�9�?l-����l��;���=w�C��i�(����>��3�ψY���r��A&�����-�0p��ҖٿL`{��/��Mlҋ�j+9r,P�Y�I&n�����!y^��H���¹`*��1]�̐�c�bqh,���5�*�ogͪ٠�?��ե^�M� �B���������hC�c��0i��Fo\F�3���lk�d���,_-���*�}w���]7`�v
���m�XuFu&ʿ�5�;�4���2���*V��h�����۸�<ݥeN��o��֪6����gC�\�i� �!Zx�ۊP8·;{֭����|��)/��6pa?9�yG���n�5uI���f�3��,{.煎[q4iHi2���B��@(�6�6պ�'����1b������w�0�S̻�M������Y�Y!{�q��R�A���)���=�p��l��f[�]=�}�B$�t![�����HK���ne��[���㋱ƣ7�o7�351�w��O04q1=z#���ُIM��zQ^pa�V��o��-2L�Y�A��/gT(�:�DV��
	�d�2}��-O,� �&K5�B�_kȼ�clW��tA(�h���kW	��ڽjk���̲C���Gx�W�GP^�p�_���\��dk^e-*D�����?�.5� 3����X���R{��{����i�& � bhC�ec�杽.�kn� �t�{C����>S�{�X�Q�;,�8e�Ǡu�!�^;��`����oO^
����)9'�-��r���]���3S�ŏ0�uhhGm���Գ�ud�)dio=a����bGL扬�+��E��m�H��#�Y�387:����y�m�9Xx���a1���Q��;I�ռ�"
#~����M\Xɀ疊EBt����p~��'#�4`�u91����Ѓ�X�?Ѕ�S����z�lyO�M&��W5O�"�\��E�Y<�׽!�呝����s5��}��!��3"���x���������8���`N�^�5B1@'k_9nkTD��u�Od`+�A�Ǌ�Cf��X���3�cH�S<�G��a����On3�th
�A��̹����sӏ�z��I;����}����h:y�K�y'�!�:���Mf�,����5��!Xy���{C����~c�xsΈ��{�F�]�U?��kW^yn��!�V�����vA�����j#}��ب�n�cL�nO~��$WI�m�w�ߞ�VPF'�tfSnA%�8�+��?���|�4X������2,���!,i�$���Q`�����œ����v�}�8��Dg���a־�&y�ZNNӅ���=��A���-z������|�- fbT�=u&:�^�;�y)��d_f�C�.�57�!�J���f�4��gT��Ґ� ��^�3�_WX}�%�|�4Y�4�E�KHM�|�^����eb�
����:U�c��� ���D��Z���Y�)��}�U��,�O�IF+U$S����;�W�h0O��f���K���w�L��ắ������"�?(��:S��,ap@�G�"A������ru�Q'���r!L���f���F3.���s�I��%�<�~,Ş�vgF��I��?���3�"T@���SȑB�7���i�,��o#�g��+0J��{Ċ��*�Z�>��5��4���(�m�*�l��ҽf���R�ff�ōU=�$Q��خ�?D�A�\���A���8gX�]2���^�/��Aց6쭑5pY
��8H,#kIo��2_}���A �
��T�~�E�nU���ņ�!B��K�E=˅A����S
�`E`�1!tH����&��d�0��Ó�M��o�W�*�.]w����عe�Mn��rGt#��[b��L����ϐ�I��RD��������h�o���y�|=�K�5^�GJ��o#F�lIQ��w�L�Zy�| ��8䶘���|e����$i��Mٸ�b�k�>�ݢ#Ҭ�鼕� 3RS�G����d8䆓�$�9��xɝW�#�DEG�y��_D�� ���]a%�r�����䮤����"������]��Jܑ��*
rM��o��z�]	�Y��,�'k������即"8A�NɬO��0֯�:����؂т:e{���G}�<HL?-ߺtĮ~�[��Kޒs�)��e���c/�V3u-��4q{R��h�������U^���Qo�����Ȏ��7-ڵ8Ե��ʖ
Lj�"��Q	��ޘ�4E*���F�1�4�M���u��B��o�����$�	8����/l�=]�!�/�<�o�/�<�ɘ��}��n��,�zB�x��v��53ri> @�quh����p���^Ҍ#��p���s�f��/3+�%�����m�_���m�g㗅וWHdM�X����CKw8�^l��@���1�j��o����Z��X"/�Ÿ�Փ���?�Ŏ��	=�L�v�7���]����[t�!��!ɐ&����,'�����ĐgEH/�ڦ�O�(zp~@���L�4����Q�؉��~&���p��+�{�@Ȉif�F�
�lll���Q��B��W����(~�5_��o���WzYC��B�8r� i< ����n��dss�`��D��_�,&>��vv)��&^��T9����ى��v�lk5��9�P������d_�_��H�~6��$��P���J<��@R�{���n7����� �w� �Ԇ�5�a8	I'Ԓ�bK��6b,�F���]nDԉt��*n��C*��9�0�z���B��[q�Y8��;!>$�m�)I�~ڼ����Mf0�i4���7	������n�E#�������=pJ�$��jlP�C�<�e1�d�;��\=��s{�H	)�ql�X}d�	S>8Z�Q���
xwJ9C9�^���7���@Ŋ��*�̏��-e��y�^��SC�۔�4_b���� ��,�g�O��;�5[I�����⢸ʌS�c�Jjis���Y�4�#����i���c*� ��R���e9X#v�d���v2�E���!ˏ�ɬ�;�����L��u�	���œ�Uu$7�i������M�z!L�@��ߵJ܀%?Mt��]?��(���T�Ws3D����E[;!�����s��Iv�������~@���ߨ�sF�sd�_9�Sj	�U�7a�M5/�ō�1���Ėh���ݕ���V��G��kx�7��� �@�oՋ�N�y������b	�䄌�`zmQ����t!��-�՛��e,q|M��L���B�3Ps�1��ũ$d%2kr��A6��2A��>¿U�v��Ы��u�*��&��x�6B�.�K�U�E������T�y�!��$� !�z? ��"��;snt�7H���\�Kf�=��N�z����Э�"KjmF癔cF���/w�վ�_�91:�R�4�haf���y�����ݕH��%��b�*�|�W����VF������V�az�j=uEI��a�?�cû��(��Ε��|�����\�'��7Z�/m��8��Z�v^A�װ�3�bϊB�P_�@��<���מ��*�D�����Җ�dIŝ�m-\;y��<�W��
�2��T#��g@�E�tC�O@{�izr�P�̏)rő�4�j;�+�)��Zov���m>��D��^{��c�ysYx��b b>?��>�`�;����<��0�U	X60	;���QQ�dR���-��
E��'�"�y�����E�_EWl֥iX
���eV�����ֻ��8����4��$#�e6� �#�+Q#F�)I:ڑg(���"=�Փ�� c�b$+�~9Y��� 
gr��k�?ܗZt������1h>bd��˽���r)��}����$M=���gd�����^�: 匨����m�;�3(��³�ɺq�>۪I�|5��$Ȩ�,Kq{8v6�X��̢�Rt~.������z����^)T��33�K��y���%�(b�n�F��\3e<Y���aF5	�.��rAwR���Z@�����"E1���M��E���E����6.�Iɇ{*�Z�<a41�'f4�:"q��!R֋��7��G�d[I%��w�=\�T���ڔ�@D:��	[�x��1
��Q�fJ����`��V'Dƛe�u������Δ�o3ߨ,�u~�u�6�;}��ˑ	8V��Q�5�m�?5���e���h��n,��X��m���>�{�\U�+\b��.��*�4� ���Ս'*��aDo�Ǭ��Wݡ�+��k���������(�Ǌ���IL�)�G��6���fq���-�@��3�C�|�4�H����b�4��!7��g�F�DL�$֮���uF.c�*�A�b�1R��(�o�����'����jJё�>kF)NP��]4��IK:򤛔>�K[�U��4S��zrN�6���9����è�z���g��ȈHT�a�v���i"Bc��TKV;�Z�����mڌ%� �Z�:ֻ_�7�S����� %�~�p+���-��Q��٦�L<r�h��K����[{LQ�E�O�տ��,@�z�j!}�w��ɑ���._�0�2�ǈB���w�SxP���mH�,A���'���Cnl��������{8!�M��3�Ӷ>�?��{�$�%�mS�V}�w�U���PI�<���� �r�ѡd"ɩ�d��N"<,_�{�z�g��&���ow�=d�Mʞ���?1꬯�:H~?�^�0w$�x둖�>��(�v�Y&��ZH8�bC�p�ż�N��^�O�;(����®�qP~��*||]�`��E��3r�c��m'�:�?=9a��Ԟ����B{�)�؛�����%�љ�tU#z���Ϡ��T�e�c�kqŊZ� 5�*�[ĸ�X��z5��C���i}Juo���n��y�$�^�":b@+Qު�ο}� |�1��������8�����B���Q�ֲ{�C��Z^i���;�C��/�.����h3a��$�>��l��wMmyf�r(O���:>�#l�o(ܰ�P�ikI©5�2 qZ�ZV���]��Y�E�n���Ɲ�M&[�Tk���w�\�X]��rTh6F`�{!^{P6�d�ꢠqG4��3�w���ƁH_���:]��7C#�G���x��T-H�r�M�q8���~��A��8]hW��2�3����1Q�Ƴ�m�Ưucs>R>Gd�/h�O��ݛ��:{�rO.���#(ѕ�0�#�K������Z��zU�-���ԤI��q��F�8�GҢ�d�����)F��[I#%+�xI}9�u��"{8J�_61��4.]\��v��vh+������f�qa��'sڰ~�*��U0�q���WcE��¡�� ZA�(�U� .'�����o+6T{7&[l���֟�.O�nQӑ��O�eo��<_���u�Teg4%��B��/�xoj�ա���k(a�j7�bY��)=n��v�E]�������;���Qy��7�9�
�l[?�k�@�:���#��ʬ�|x����������*������vo�V�Y}��4�`9UG
��b�sK�X�"Bp�a��d䨰�]���Hp��Hx��N�6>��sѩ���,��"���)�[���D#>4G��Q�=���;���^|�s]�I�o�Ώ�nX�f��&H��5dR 8v����YJ��	�B�Aҵ{G��1:�+g}|�<1b���PB�x/�b�k\x
�0�
����ٽf�}j�����$|�>[�'�=�� ڣ���o��K���V��z��/Sx����4���mG�-�+���F�]; �Cix�����8T�B�� E?�H'R��$%�����?-ed��V+���+p�5X�G��o������������*�lTb��O��X�@�+�Rnמu����]r����x��8tc��dş�FIi��)���/���a���L��1�8�f<�U�C����d�Ρ�J̮:�~�E�)�_{>��X��'9�;��h�9-Jd���%�L3������e��!\��\S�x�:Ȏ��4&��X��<0�D v���{ܴ��og4�-�g��H�2��5����u`6�$j�h�4&�#8����(�PEv�[�Q|5q$��9#u�V��=���Ε��7�9�\W*潌A���NE��̷���e�X�pk�Y��&�M�Θ>!m�(�á�ȯ�	F�M��4�y��dI�`����ϏD胫�gRO��p�R�p�#�����=��d@Q�ɐWK;i9�=q/�q�lC�:�ޞc�m�>w��E���2���{`���`�R��8paDIϤ�^�9��N�r��z7h�]��٧���E�u����4z��W�TZ�K�L|�K1?�I	d�׼UJ��e�����������W�#��I|gt�u�"�ׂ�`;��(W�xƿ�s�� �%�gp����=>/�Mc����Wo�d?g�
+cg6�QB�<����� �ն�끿U着W\.�_s�$yK<Ȏ`� ��mS�f�V+��`��QuӶ�VY��Gʘe[��9V|�__^o�J�
x*_�֬��vt�fF����p��N��z���\��nO�fo��Z�����e��mbPX�q"�n�gB<�\���Fq��c��æW'}��9E�7ǟ�R@�uX=�J��N�<���UK��IX
b���Ɩ��C�}[�=�/G���@��Xb����2x�Z!��+����ף�-���H���~5(�˧߂9e�IjjdYI�^n+�����lk�V⧅���?��Ӡ��1U��dHO�E��
o��.�a������.���Zβۗ�hzp��p�e��n�
@XApps荠���H!��,�e�_p6o�ծx[��x ��I��ۓ�|��ֿ{�ZO��<M�IG�1����O�}o�9�lZ�� *���3�����`�^Ei�������%�-��yU�;G@�#�t1i�0x[\TVh�[3v���)�pYA1��n���󢏮�P�|+u�L���|5�f�t_��������;�ԟ��u5	Q��┪���Jߎ}��_Y]�><���Ro�NX��)�گ��a��e�M�\��R1�3�r�o���+�{ fH��Q�8���ui�G��mH���x8�I�_�]��`t��X�N&j���"}{+|Ϣ��R	h�vw�f���k覧8'h���g��d�#���'���:�e���i�3�[��&�۴�;���r�/a�8)	 ��S�|تi���w?_�(�=Z���S��]���G��#�ǻRDLk��J�(.�	ǃ~G�$��.�r�g�fkR�*������܄�s8َt��za�O���� E�c#)�NE$�����7zݪ(v�)۝K�c�b��Ȭ&[���	S+�Fʻ�Oc��>Y��G��xNe�sUN��dfkqѧ������7nOK�R��QW��Y�
��1����纨̻��a���Ӄ�#�B�?���z�Ք��4P���T��L�y�!�����}�e�X���͙��N�>�q�3�^�
}�SK��n�� MfX�B�E��"(��Q�R�_���+o��y�KQ���8}��m�5�,N>�?�
҇��!h�t��mTٱLZ�K��b�9<ds�_��j�3�$��C�o���1xՉ����]P�v��u��}=}�h_������]�кR�3ut�&�r�����B���`^��)=�gƞ��E^)�C^bߥ��!��̎w*`$��)r�27�憊S�����s8/ID��k��}�7G)'�	�>�K��D*�{��TW��n1���k��z��ym�vI��]ٌ�=<���Q� �IQ��{j|L,������yt����b͝�)��t�p�hbl�Ƨr-��	�<Uw�V��]Xy�΍7�K��������+s���;�;�B'[�s�8��D@_���Х�qxak�������κ���Y5�u��������V�$qƍ����a�^F�~��݄�E��'�l
���Ԉ��
9��z@����k��c����;�o�	x<��"�����s!f�����$�^���[p=����Y�q�:�κ�3�>��
O��@��zGy\ԅ�������i ���8�,�S P��5�\;����Ŗ:�La�/'f�#B�R0��7Y�ϖ��-@�2��;V'��$/��h¶o$s��e��:j�H��M�D �j��E�M��j�@�0��'_5�T�������G��8«�Љ�Ռ?� ���~��W��F��pq¯�.n�8I�jU�Bj�H}'TC7�3<����u�h2���з��CR�':��S�S�sRqzt��[Ii�� K�$������� ��t�\��E���������ߔ)�����:Cf
  7��5� ��0��u8I� ��_z�2Q���i��z;�����h�d4�u ��>\�;#F����o���,��kp��G#ތ\PVm��v�fQ�q0��vЧܭ�݊U�N@.��75o7�J�@��L�5�vi�i�`�*Ɓ�����x�N��N��u���N�>��`�2��=�	�j�)q���>�A��m��r)z�F��<W5��[	�~�v|�V>!��A�'���� ���*�a��ĥ�Z��A�ܖ>��U��ܑ�uO�s�(+H(��GM3����R�\��ORa�'>���v�9��:��l�y4�d3U�%Zߑ����A@���Z��&�F'��N��@���7˚)�wU�-�w�]/{[ͭr_�m�u@��Fѱ%�QKU�&U������eM���c]�$d6�h&�వ S$1~Ԅ ���*�"*)]b�Ͼ�U@k�2�+�6Nn5d�����F�k^�%�](q��.σ�YF��QD�.�2{����i�%5����;]�1	k�*6n,�˙�a:6����c�	;�@D��4�}��,��;�����+��4�zy��Rv{Ȱ�h����I�>%�V�CL� �9��4�Li$�l��j��-���x'C�YQlF� �J��[�n�y�����E�����y��PO�۷�����W3˕�꩖D�UM�����L:C��\J!(mFg:|��P�Eg��oqױ!n���n����!*&���'��6��� �S�:����PǤ��XX8Ц��Kz9K�c�d*�J���{V$�Q�y��Gx��>�|3P�:s+X�3;0R���1�{��u���ӡ��B��,>�M�o�ܼ?G��R|�#��{SI��bhS�ꭆ�i'��?�bQ� 6F��N݅إ���4|��5��H����V�4\P��e�9�u�L�$�)��w��wY3�7Phma�A� �XH2��}H Qg,��6�~��q�5��P7'���4��O���)�YᆤtB1����~ܽXcC�h֭��^I����gm��N��ŷ�*����"@�?J�҈XF>�k�Èx%�u�C~�2�$|�0�[����W'�se����&v�"�����M�=["`�i�M����nm��Y�6��-�4�D^h_�"���6��jUq�aGE8:ʨc`v����C�I����5��QD� �w�J��nO�Sٗ��(m��M�V�P����:9���D�ק�6�Kp���o�/����O������_�BDݹ0��K�˫�7�;�E����jr���i�B5�C�{�w�$Eм�2\��{#���;]^�oäɯ7��n�R�� �@� ,ͥ2���ϥB�&����܍���$��?�Y�ӫb��_�6Z����<!��q�����-��LGc6{�P��{��|	���Dl	�tL5�$p}U0�G���������t�x��X�dT�}|ӏ�Tz��PjDr��ں[9mҝz�K��hj�;�}O38C�l`3lJ�_)�-Z����핲(�J��Y�W�d1|�GG�6��J��;,���~������~ɉ�m�L�.b"�q�Dq�ѝ*�fBe@w9�DQ]b�|����N�K��t~��cI�Mb�K���^pF3"��Q���P�pf%a7�n��?X��<e��r4��rSf8�Ұ��Mj:٭K�y���v,�t���
n��	�6���'�A����E}�T�4��k��s��f�l>{�T��M� 8�'���Yx˙������(� ��9�!5��w/?jI%��uG|��{$KX�#/�8�fqɿ,�!�Ѻ���A��Y�9~����=&Q���{�M��E2|�fT�符��@�������[��o]�M�"r��t�Y"���ى�isx��[ 1y�)�76�9�{[¶�u���1!�Mr��4����Fኝ\e?}��V�V8!YZ���mA���'\���	�ib�{���ތ��,��-�z��Ō)�N#h��蟿4W[MX�]b[��ͩ1�����s�k��P�˼]-��Өa2"b��$ ����7�8��J�9I��ʕm����+3cմj��*t"tK�aH��`���"
h"�:Za��;~.kͮ�f v�pb6��򽦘�+���	X���d^b!>�\�s�������I�o`�C���W�%'��
<���D*3TL  3LbF�1K�Ũa 䢃G�(S�n\F�j=����9��Y��dr-T�"��V�d���b'�(�������/���r]ܦ��$E#Z�,7��ΆF5;
���}����M�#��������a��
�$�V��'l��#=��;u����qH8�Mbpt$����}��&�1K�U�/�{��c��E���S��v��,��VtW2��)Z�.���=���ZU�n�w�掋uh1ʌ��H�E\K~�΃Fv�Jc
U�.��A��:B�y\��!���P۽ME]��J�h&Av��׀�8���DUm�iZ
ښ�g�J��dk�p�Cxqq��:��86wՐ�(��|���z����S�j�@�|����z�W�-mƲG������p�ɒ�sm1�&PD�c���BD�!>E������x��qk��T���'��'R ����*,
>���]�
o/蠾���L�x<c�>m���.� ������;�s�K��(���H�
���A�Dמ���N4Լ�����`B7�a���b�e��-�K����w*�eOț3��i��C�%B�<�K��Z���;�v^��B\�I:��\��y�UY�K�)[�r-�E��%�Z�,�Ǉ�h�3�0�Z���1n6�󟴗97V��R���{j����H��.p~�]�K����J��su�dmr�L�=TuBT+�����:w>Z�D�3"˜��E���/�Vo\uU�%0���gb� �)S��ZA۱��yMe��iP���z��}dC�P�(�xԗ�[��FQ�d��Y�rVDu[O~*���b
�GƟ̳��� .�^�&��ڌd#7����rU�:6�H߸*9/|�
i[2�{�~���m�йZ���V���oL�'�ȵ4 ��V��B����Vre���U�l�S�]�s�E
���2&��~�Ȇ	5�d�+e�v���e*���o,���3°B��n܊����f��TX�7��XܘCD�{٪\��)v������-����n��T J�eQ�Z�ϮrU���2v/$��U�$3����a��b3��M5 �$#EMa��|�NX��'���c�g؉b��&�I��Wl�?¤�Y�ޒ�����*�fm����*@���(n���GLfj�[��[���0D�Ĉ����8g�����������t�����ӳ�)���)͒�c�瑼����K�p"���������ZjJ��ߕ���*�2_Z9tlfgT�8��'$�g�Mӎ����L��yBF����
����	)��,<�n�A伇i�E�?c�N5IQ�ie���4�Q$��7�'|2���@S�(e�Lr���]��;�oz��-��&Ǜ��]ǫ��n�p~������R���E����]�j��>1Z�f/�'=,I�!a��v�K�1������]�{���̥rY����R? ��Zii�̐���K];�ߊ�w��Zk�(3V�^>������7�r�yFD��5��A\�VAr����`H6�f�����⪍�.p����$�&��qf���bHֽ����,7^�r\�_����	�<��iGQ��&Mﲬ�׸�S)��@�]����g�����2륺�q���o�ҮقDU�-reQ*
#v����=6 ���?f"��+��HUX���D�C&��m?�u�G�1͊���'�A{�f���A�bk�{��i.�ct��_4�bStj��+H��4pŅvɿ�1��+����7$��U~����e���:�i�~�e�Ba�ya��W�7qA|&@O"�0��%�N���c��e]�0���t��(�^�Y=^x[8=�W� M<�`��K�U! ��<+yT�59��v�91]��e~������2�=[�2j�Jđ(�,�R%���J�YSucO��Z�~�r���[wRUPR�)�������&���������ɃKz{�bFA=������D�TR}C�Z4��рv�yj�G�H�{ڽ)>����}�25��4�{@I�zQP�1�������8�G5��N�h,4ٱ`���en(*����{
殿�Q����Զ�tU"���C��QE��!�[t�1N]�I
B�e,.�Xq�V:m4{#wfcpRe릛XF�4؁x�h�z^XS#�7X�MP2�Xx� ��A��!��K}�� �qp]()�����z���A�����o�5<~oN�%c��#���|m�����5��r� o!�V"U�[:{6������Z�9�ǹXK�3������fɁfn�ݮ���F~�n\��_�O�R���B�o��?X�̻���:��)C���mHU�;\��2q����wKj �ɨŭ/Ev��-A~����g�$��.�Y�9��f�곀�ֈ�Έ܆�xg4��[q�`�a����N� pSNǟ��E�J|(�-�zr5�Z̊����Y���M표���Y�n�p)$�9�˷���7�~sQ:������*1V`Y���	�B��B���Q�;yv��Ew�y+��3F�f���D��-�7�_��a�2e�1�6=�ΰ=�������h݃ݵkkpQ��'r�N�b���⹙~�):�:�z�+U�,�WQ�`�M�ub<���.��������hD�݋[�ѩ	9i<)Ħѥ�B�4<`�mQ��Ȗ�R��dɊ��'�`����2z��Q��~��NWq�����	�&�٘�t��t	�N8�Xi� ,s�B��I�]���R!#�}B0��#���nz�?8��a���ԭ�D55#ꮒ��P'�^����H�`Hϱ������5�vvrC�M*A�����3�9l�:��?���X��1��h�7u��&L5y�k.�V����V�� �8R:	H��Kr`��W�	[��i�_��b�����l���L�����{6��vΥ�ʓ͝�NyM~������Qf���|���MƳ���;�plX��Xa�l�MnCp�;����9S�Ъ�3i�GTe��U����f�*���Lk�s�{F\p�_�	6������2��r���.�/��sbn���Mֿ�)H#�![�
*>�1������ G�%���������[��Ϻ�?)H?�B��b>�J"/�	pL͔懶���x�e�>��᷿Ψ��E������`���f��-�4H��%��f�<<^����R5Z��HX�;ք�h˱�+�����ó�݇�r� ���s��KC�/י�uC�Q^��5�}��o�R��۸�������N�H����cj~���.����)�uz��y rI��$���,���5"��z����[�Dךm�2�\���S���I.p�[_!6<��[�P`��6F�Ѩ ��-�G��ޑ�����qb1�7hJ�a�?	V��.��8L!q���X۹,:��\����nK=��u5|�٧	{RcI�b�Ϲ����2�.QC^��6�}eq�a����;��3�-Ϙ�9�%�Ӓq��h�zK��w��D%��"�7�$I�Nw�W�𥧉jV�Q4���:ш���^9W-��-LK�W�\ឞ��K���W�"�$B�J�7"�|�^}�i�|�o���,�)������q�<�S{�F�����.���1����a��w���^�ݐ�E�m����{�9�B�2�_7!������(��A�8dލ�kOn�b�X?��PUKQ�RWl���K�vcO��dS�@�Bx��r"ڶ��ΠV����J2�Χ?�9�wnk2Z��^����?��xz�۪8�P���E�:��Wk��޵��JC-"����t[]2��xV���F��w:b�20�~oյ�l"���	�o��"� �I�����Xɥ�+�Icc�Dv�%$H�<}\gU|vB彤W5@ƈ�b�?N�$���q��#(��(R#��!�Hʣkx�-��]'�.ҋ�;�s�"&@��]�0�V��G
p��k�m[E�W����IRLbDȧ£G��V�D�/x��-�7�����/b��2�1AzJ#,�2�9Um���1f�f���<e����	�^m�{b�[C\��+��M�� �I� �¯0�Xd7(�ؒ�2��JH{ 7}�p_:�M�5SP6�I��ЮD�e=2�M��g&=N��Q ��s.D[#�����*n�cu.�X��?s�<W��A�j��h�^x��+~6��!�\�%��͟����_�&5-]�3�w��H4��b~�֗���?��{g��-���G��$�[���0�ɧ_bM�A}�h��1{���=�`�	�i�*(�A��Y{jP�A�"#x����Q���}�<��GM�F!�?�M�4��I9)jі
q4��f�,�3����!Y���o��Hf4�l�U��l�/"���@��3S��n��1���(/�`^�i�yG9{ �+/wsq�'��Mw��[� &Y�h�,�tz�j3=|nN-��a�A~�o"
�@"Vo�9�k���:�:�_Pٽto�_�q4�5�"g��nX�S\�A��� <9���l�X��y]|�׵�G;�O���Th,�����_��lPs����Zm�~叧�:�$
Ё�1�������C])ݧ� }�E����Ҭ�t�EG�qs'�`��+�
����j������Y�c�;�*��Q8�½�^�����i�Ott�zB�6?��Z�Ô1)�#6Ui}М=�袒�g�/΃ -���#x2�Ib1ǹ�h?껀R�:A�'@\�Yj2A��'��	�kΑ5¨J�
� �������(R�U�(Ea�`�DJ��pnv�ť����<8s�ԍ��==>XN��J���ӥo#�@�7���H,<��kg�@�& p.���%��_I��gQ���M������΋_|^�l�p��XTps_��Ͷc�#��ݤAf��P4�X��W+��yݛ���9|#�dqw�k����/�́{G�m��Gy�`"}4t���`�ے0�2b�ܯ܈��r"��[�l
��O��Y��@z��=�>m��y]��r��Ȭޢ�Z]ve/��)�psgRɸ,�t�U~��	�]�İ��"s�q3R蛖Oe.��6�*}˶S@��lS ��$��|Մ� VT���&�F{�v�~Dޒ��v�uN��˵���\C�l���J�u�P�Gj�`�K�|�K�K�g��л價1��c��8TY��m=�cY��WK��ه5�<E^Cc�+��&Ђ��1��@d�s��0������.�^��x�g���䙝vN;�P�5S���ި��£C�9}3�L�s4��(.��A�azh�Q��R��G�KqAT9���{���-<;Kb��<��hq���V�`}L����sO�Y���g�L1~-����a�D�W�_�m�{5�N����_^)�k!��~ր4��wFHJ�m0i^�ƁS�}�>����o�UR4�Q�á�v���&1sg�"WX��ҷ�@��{\uH4$c '�vjՂ+�����6J�pI��/�+��+ЕUrc��7K�	Y�<�{9V�b�+ܨ:n��n!s~���U1�e�9Ā7r�"Im����+$h���^���ʋe�o�BJw�쭴**ư�Ua	��Ң�N����o��J�L�_�5 �1��K��zE�:����<M�,�.܈
ߚ�@µp%x;���)�U�a�7���s�,6l�#<�D�~FbnM�d��~��!ڐ�*���9�gt���j�����HgdCW����yd�KT�j�{�Ru�|�Q߼�2h�e�*g	�Ln���?�$�;���DtTgZg��M����A�9F�';�]�-ݤ��|����g\���^z*|�'>Y�׵��s9���[T�3+�s�>�b�Л�����dŲ��@��-�ot��K��������
V{���a�2����Gt��ߌ�폺����Qu���*��<ɻ�g�5Ҹ9-��+9�.RIǎ�)�9y��Ub�P��K���Y��;swջ4���(Y�ݗ��z���4��G���M|�H�ab�D�,z�b�����~�[�ީ��I�E���K������"����@�RqG �:ܢ��d^+��{�0����vg����EM�!�9�	��O�A��at�R&�Mꆽ����(/��Xc������2�� �$cB P?�V��5�@��r-Cp5eH��,�i�,gV���uD���Y���v0���.��a��}7w��\%�k��Eܨp�"�������"� ���FK#"�ɪQՇ�em%�;6I)Q�P��Aw���Z���=�2*�ܰ*ǉ�*����+2%P�+�r~=R�+LtR.�$r?���	�/�kV���-_�x�y}���PCY��k�[
�~FP�i���\����[�X.�6y�����+�R��'��"���K�]��Ͼ�X���4�u��D5A��.�t)*�R
�|��A�0�L吚��a��Fj�[ gܣ�+u�[4+�|��3��Y���H -�H�����<ibiE���s��޺C�L+=�̊�̎](������bx-2����%�g�$wa�Bw���	��۸h@;�X�g����9(̚m�t��T�>�9�a:9�q	��N����
N�?�24�^4Kqr�f?1��Zs�)��,������`��P��݁A�JĮ:�rQ�3�[?qZa�lN��xc���q_�"�:����`����8�>��4ooѥf��o(��܆��]z=��|�������N���&Ո!�\��K��l����=��e��wg�8Ulm�����W�����j��A9T�e�g��.=�>,�2�
t����.2�Y��B��q�X�_ث|���nB�h��=	@6i^0���9r�Q1籓I\��v*n�����W����,�����EP'
V��|�p)�o\���S��G�8�	�1:t�Y��㠼�L�5t8��*�Mi��X!��I?�+��`JyB]@Ŋk��[{�l�vX%[~�_1�?���X/�]Vuf���`&���@��A�px���4�vP������<�m�S,��F6��xW���R���O��E	=��m}�V����)�Z�����z</�R�;ړ�~~i�������/����kB�� ���i�l��G4x�`μj�D��,�M��iJ4����[��::I�څ ����*�������g�����H��h}vj�[��3���&��6	��$�����ڠ�~D؀z�N�5�����LN,A����g$�Z����Q���"o��/�<C�j)�8B�
�Qe(Ry[��@A�.}�Y#�85Ke�|��n�(R��f����bΥ��9��ҏ��ݣ�x:W����'@֙A7]�����K���P�_gr/~�O�"6�k$�2�9�����h�Y5���u_�E�i(~܈sl�=��'����-���;�Q�=��H^s�Xg���[�� $>.P]�V�Tc��fdXb�������I;!_E��'����)}�:���G[���+	�ݧ�O3��|X�(sM�0�/�׾+D��F����^S;=��^v	����k	�3H�s�a�� �͕��O�w�V��WK��|5'/l�-������Q�c�w�6t�w/�����m�QW�*��`�q��S;�۰�zS4��Y�3�H|8UK]A�GJ~=׆���P�9�Ѭ;7�;o�'�ff��<i\�[? ���ӫ���e׷}��mw�r9��=;?h^�X�?�����"�5�'��ˌ;�O�w(�K�5����Je�7���݅�b�8Ғ&4�U���t*R�:�U(�,:wm�2�F�P�ݖP�@73O�I�-��)�&���Ns�ɩ�gm�M�=1m�x@%$���5p�Vjd��ۼ��Ht�6��9�M��ƨ?�\�������.C!.�d�|�t똞��'�{cخ��L�ۇ�_�|��Q}�O�|��8�8M��"��\&��Gr�hR�߀Q^�'3Y��m�$��wrGc<u+��<?���>���(�^��H�]ӷ�a#^k.y%��M�(K�j���
��`�J��=^�a"8���*��.��nh��`l]"9����M-�γM��V�k�u%�h�vV%s:���k@���ia� ������['j
t�>n�]r�L��26�.c����r})\�)șl��x�`j�p��i�B����,��Nj_�U,q��Z�� �S�
�����x`FO�P�+��0,����h� �,5�:4ܠ��X`?��\w���.��z��܏�W��z�*w��eޔ�;���B̪9;�!]E�������W( 2�/�l�F��&����̣�ė�Q_[�����4�8a���{hBK� V�y }	iPU�m%񓇼�lC���7�$�E��4_�hQ�B��� ������o[�0a�
N�2�鼮�6���)����8{Jw�g)�Ļ�Iw����8y�E��l!�k
Y�rċ�A�j���Rqpbp��
�T�K�ٜ�#����ދ�����T���ګ/�.�DQ5���a��H�p&�zR��� K�/�&G�c@�������dP�R�?S1-Ε&8��|@w`�W���#����dے�4�d]��`O���H��`0L#(jD�q�z�]=��A�fo�vc��4�z�g����>�ı�Y4T��x*?�Be���A�����>-*��~;p���\�$=��\����|5R�66W��ZI!t�&	l�wP��D#�Z�ecs��6d�c1������!���z�s3 �ufza+fC�!����F�l"�����r�G�ܴ w�������qC��P1?�do[%�\H�k�y��k|2�诬�,� �eF`HBw�uǥ��E�����&��)R4�Ҹ"�P��麙ǽ����]>��o3{Ʈc&�C�����_��}�����]zH�����َ޽�-�UZT�$�D��� BqG�2>}5��'�Q>L��/���t������㒪�>���i5c�<S���N��rT=�� ��H��eGÊ����J�%`&Y��~v�t��"!�wz㲡o����$욙h�񢖡�A��-}�R�B|πeqy|�F��.~#p�PjSaNvo��ȋ�_9GC�r2����ؼ.R������[
5�Oʂ����ʒ�g �_%ڎO07g�2�������7��D3`��Ē{���m���KP��ê�ͦ�j�أG�#h����p����اr��R����'D�/@Ⱥ�[��y(f��࿗�v?=d��ۯ�G����'(]Ux��Iw�9"����af�I�C�"��ђ�>���J�%d����ޏ~
z��m����i�&����MAcW���s~ք=�����5Lgψ�����6�=�dRV���l^,�ɛM�=1�板H�����v~GQ�cl_�ba��k��fn]��Y �(�^�A( �S�*�+�oqO�J@-:����o�4Ŝ���x/��N�#�9Y2],�䳷�q��B&@7z�+=�_�e�з�5�x��Ӝ8��������r�VZy�C�_��H����v#V;�y�R�bU� r����k?`��74֎4�g��i�@�z�v"�If��&h�p�s�w�N9L�C�`�Q��U�3?;��o�&��ƞn���+v����dh9�(���E��AJ�U��M�',�A�ޕ�5|�z��Z߰�� �D�P���:�ӂ�8�a\O�6js�̚9Сu�ث�S*!G��>���LK����eG�6Ck)P�:�v&vt��J��_;B�j�P7�Y*�p;���h!3�t�ɉc�D��5A���ޣ���A�I��_��b��l"�����ѮT�b�+t�a\���%P�٢1ץ�-w+��l�
Usw��>sOƉò�dρ��������\���ś�]cX<r��U����&9*�rw����тS�EL�W�XvEIo7�������2	޸;�<�pXIzD{�ϴ��i"��|ɪ�fu����:Y��/���i�A��`B��{َ���<D�
�;�F��)g!��7H@��p;ʶ����
�q�]1���v�j�����JO�y�a��R����{��	�R��H�W�k���YD�# �3�%J�2_�{G�
��e�o�A��S�ه� ��)2�P��y�{�L}� �D5!nW/U�u\��(��I���������)'t��>����h�G�u�sh<#t���\�g�����lt���vv(tt�w%]�Z�V7�iSd�ϴ��A n�}II᫊4�5���MV�d77��f}|2��L[�I����F8���Ԛ+S�`gZ�Gx*Ĕ�����w��͘D.��D���|# Mb�;E�DQ����i���r;��Z�<w��q�#z鶎�mPi]+@0OJ�S] +7R�;���x�=�))�$Ng�Դ	���͠���{�Mץ���p�����A��t&T�m�����6e�#+� �#Da���Ї�a�7LIKK��lVh+�����٬�x�g:<`�)魋��Ӑ�ɍ���d��@Ե0�{���`�u3��"ҍ�0w���������vA1�q��[������@+a��w�96ŅB~\'��ˑ�<9��K���d�i�U�7�^�~��H;Kgk����JQ�����u!��^����v&�]�>T>_�iv,��g����ͅf�uտ��w[�7|N�$7��JD�r@���g�G�5�w���x�QY|��,�*���Np;�ߐ���`�wciE}��B'B��^U�"ʪ[�ۚ89�̝��@���n���۹e�t��8��S�6AKD7u���b�A�9�ˇ�xl�8'R׺8,u��T���O�;�:7�<4	��XD\V��V�s ;lJ���8F"=��r�n�p呃�q,���%�����e�	�ib^�����Q#��ίM��~��1�87��(_�qв��bx��������ybqQ��«�iM���@�n��z^���S�����ӣy �(ȇ���\WY��)<o���"�}iV���� C�s&���~P�m��:f8Vdj���C�u�M[�(�?+�Go�����z�����^3h
b�v1�����G�ɽ���Q�`,?���3(�'3��@a��Rh�蔿;ǽ�N���`��7�g����ha'���IQ�[�������z���OI&����}��l�Т\S��gq��0�i�)7CP�*�H>����ݦo6�`^����\P�B�A�
<#>��"柁���k�[�_�)�ǂ!c�����S2���4�О��v�T;kˑgE+���
J~TV<2_��������H���v���fGgt����_~�2;r�p\>R�D��k�Ag�=���C�r��5���>�p�#��!�ܖ����
�`�s������媜z���?���ϱ�$�c.s-���κ���O�$�� 0^��Rŏ�(����t�|H�/��㗽D�]�xMF�{/{x����䜥Q����i��?٬
{�Ey�1*�ӏH�9u㫤�F�"2���0D�o7GT�N'P�Al�	D��W
���	����J]�	�Ҫ������Oowfʪ�9=~&࢏�j^��ܗ��K}mݛC�,ثf�L{���b��Vb��` ʇj��v�
d="5�R�[�!�F[��:�Iv�Ҳ2�	�,���xCD�����mިB�gz�6�5�ﭢBå�eX?>��S>O�n�j�3���q�,��+`�7����Eҽu<��� �/��X4\�`U\x�blLZ�zDqz=Q��돺�����3��� ��D��o�iC..��:���}���ԣ{������7"���
R�0c���4��=S�qґ�� �u��S�C�����)p�=k��Y���m�������b��kt��+r�E��MqL@�VT1��lY�9��y	Ń���R-h��5?�h�g��l �J~����gP�	孨cS@,�b#Ay�>��;}��Z}���"KLp�0�O-�vlF]e���ָQm�\��t�z;IS^5�R�tG����-���e�k���
dd =v�� -+�����~������0����؄��	"`�(���?��P�ZX���@�#��:��C�.3 f>O
|��,�S���J�Y���5�-��Č$`�[�LZ�;�#w���bm�c�����\�n��31�� �g�C�ނk&h�*9mO��T�ɺ�������,"�9s�����L,��0��^�����ɝ�79ئu���]ɛk�^���Ъì��"!��JkGΚN��U<����~��(Fp,��z ݴ�L5��N������l[�p�ܧ����>o6woo�E]���q�d1��c�F��?�%�[��!���+���|'AQ<�ʫ�ֆ�/D����F��i��W�V��sC�i�ԸV2P)�xQ1��F�pg�z^Lc��z��4O&�CW|�TXܬ���l	�S������A2��m�S3�v�wx�Y�.�R��Tg_�z��:�x'��8+*���6� uU�_?����������A�W���uB��h�r`��;-r�;$ ����u�y�����4z���j���ˉ�#ʌ�Q�}8���I�V�� "p[S#=�#_Zk�8ߴ�ԓ��P<�Rs�k���O�FP�~��zܦ��6����8��Bim��.����gg!}��� �Y��؆%H𞴎N�54�R��8`r���h6�|Y\���
�'��W�?���;��!g��0'M>�|Q�s&u�̓��_���T���`p5tվ��n�M�ZW�N�F�DԬ@��lп\��S�J{UH�f/��Z�{��o�t�oC.F؍��Ή���h"Xח6Y��J)K�c��k��P��T��ܤ��/I�*��bs�x��q��7 ���M!�t�,��th�E&p�_��z2P7K�l�`Ȗ��Bۘ��p��}�Yyy� S�\����`�پU��ؐL�wH}�Tu@qTğW�]7
B���=�2���UmAĽ�>/���0N)���pi��0���y�?@�<G����I�����"�e����F/�?����}e�m�&�
�b���^��C�êh�
 fs�VU�WC��������2\���K��O94)��h��Q	�Wi�K�X"�8��| %إXG�tb�1�Xq�iW��*L���O[A��v�pgs���`yag���*���	 T�*>=�<�h _��l����6�^ͮ:��0-��s�Nli5@>��G���d���"�"-w��QG��f���D�1F^�1Qmk�������kU����:6ֱ4h.�-����~ַ4�	(��k�GDwg%�O!��C�4f\�Q��+�Z�By�.>'����,�:^��c2�Ʀy���u���b"7W�����e������3��c�\����U#�(��i����\{�C��<l��XQ����~*��e��:�y�<�=�9���BP!��֥v��;iD4E��m�Ȝ�ɥs֡�c�zy�ǽ�(H��.C�F� \�����7���Ϟl{uM���\ ,��-�q�"��[cfQ|mO��PW��=y�p�k���B�|���^�rD�"���Do������n�om�%?�n-sq���̉dM6*�'?C�A�__��f�o�*�7A6Ɍ,@#{�K���;18���Q���Sk7VH��p{;��q��¨uA�F�z{�mj�ë#R.8�j�J��+f����4>iǁ��Q2�����a���F|@b$\o��hu��N6�Ŕ�M�Aa	J抲	���t>��UG����{ٶ�l�
�@�L�Uz���|�[�h�e5`SUq��5�z��+�����!<%v�:0c���6�7hyy�u�1D
p�]�d���{#\�&%�Z�<������>��A���ȀN�;.o�_E�
�ڑX�e7�Bh����*�@��S��|Ix��zh< ����{�[��u����a�
6��"���k�8 ������ �=tf#Dݠ�[��4�8(�F7���?F\=��Rh�=�{�El�w~|J'�ʝ�d���u\~�Ul�##�E��w�jș����r� ��:<4[u 
fcO�jgİ�\~
H@U�RM�|[,s�8���8����=D�Ũ V\��s���k���:m��W{<8���<�H�gı%�Y�(��PUc����S9_�w ��tF1���-iи"��%��U��{�I*��+��>�?.'�d�gy�,רP�5x���/��aRO����^����	��|Zu�("80m�%ͦ��*��5p�N��k�J��'��X+3�T<TtF�Gv�V��Dg�0��L11_[�25l����ձR@^��G�(���oG�Ђ�S+�,��Q�J��N
�W�5x`dO��<���6[�zt��L�&���$�0��]} �s�{���{0�	��"���_���_�܀k؊zuy���M௉u"bJ���	 ��6��C`a�Wz�{m�������e�hk�(���G����5|���-�w�� ��$)��bP+F_���"�FW�#x���N=Nl�}�5�_��@"Y(�be��N�J�C�ѻ���Bx�Y���(]_���+_�<K^���̇���0/ڄp�����@��R��_��v��r� *,�|nڣ��,�.�+HI
�0q��^,w��M�E񼙴\�=LH0�&���f{���|���1�ΐ����B�|�u��`Wy�Qa$D���d�[Pw_��1�(�uo,

���p��x�E�>G^j��%3g
��h��U�r/�Oktc�*����=1@|k��P��p� m$����-�|���d�Bz�lg5;Y�����R��b����M���5��zj������<��c�cR�~6�Gk4��W��q���\^�*�d��)(Y:%���Y�M��&~���	ҀL�͇�����I��b�'��ȯ��&�]_�X��F�O�7�lO�㞃��ә*��LX��8C������@�S�k��؊��
G�A>���~��I�����gX���\S�,�O*G�{��0G���4�'���D��v(F����ȴ�]��, L���ǬI@��Ps{��۹)Z�8�tsF� �#[�?K���J��u�YOܖ� ���٭9���gM���O�a�t�Ʋt���~[*&�	Ժw��P]��,���ނ��쳨$��@�*�t���?��T��w�W1 �R+�6<���,T�1"1��jt��pm�	�( �ȶ����-��^񦍆h^ด^���e��@tK΅����,�ξ�90�o��x-�ә�j�Y����[;�6}�ş����:���j %kJ�o0Q�OB��!���B���*���ҥR;���������h�ݑ$��
�M�P!�q�x�(Q	��f�bw;�ڃ��>��� ���`��?���������e��B����ғH�	-�!�}��)A���<�f kFV�nhH8�s��W�jF]���hn��՘ЋbkN ǆF]���c��%�S���(�j��c)!Xs��-�λЧO!\nPz<���K�	�1�
4�o�WĐS�g�qO���Th]ey��ku�&|�2��u[���{�6�ɟO��=����(�Z�O���0PW�f�3o��I^�N�ܵ�b�2c��&qH�����%����'��&��	�EKM�O�B�,��E��5�=,f����a��\BSl; Á�p��� fRhU��sDsjk��@z���a�[���Ѝ@�I�1we֢��;ZT�����H d��2,���o��4�'GQ'F�p->�!ɬzq$�P��r ���4x��*-�GA���|��1ӄ�P�,o�\4�Ӝ0�K�ͺ�n2t��s��j�%���N7��ȍ̪�>.�`��i\��.b�+��ȱ��+A1����)M]>$� �����xҺCŎ�*U��S7um�Z3e�bS�/Q��#۠�H��AR�߾7����3�pQ���b��D�N��v7][���H���[��Ɨ�D¼�X�1��#3���c���@1>B�&�bPgn��ݕZ�O���b��xc;O�#��Z�I^��g�=�������G��$���PP��ej{q�nVq\&&ܙ� ��ɀ�1QD�O��^ްy~�D���W�֧��xn}�wiLm���jȾ���xd��oLǇ�6�>8�-.ċ_�"�ey�3K59C�Zf�=mmj�c7T���_� +�,Ѩ�
�fJ�wh(���(�a����a��H���9_��Q���FTCL��z?��p���@�+��SPy�C��{��}�t�Fp�`�� �e�7���?�o��@��d}9��� =l*j�B��J~Z�cGV���Ŋ�}Y����&��s]̊�Ǔ�q+�,�����E�;{Z=I=��|
,���	��$T68LָC�|�FvG��&	e�-ul�X� Qp����-�������5$@`g� ��:K�8}Y.�{!S��J���/�6|a^9�L�Q�`�,��1���� �6 ����Y��$E���)�+ji�Қ(�N�#�bx��U�R�G��,�����>o�brP6|�S�	�-C}�mh�k���rl�|IJ��{��J�6�݃�6V��-$��h|9��|8W��-C%ƙ ��b�� �����v�ǫWTr������0F2�܉�$:��fFSy��5	D�b�����ɕ����
{���=���h�^�`�ܽ$def%�����Y��¾p��`t"�ʯ̵�^�R���C����u/�R��_������������c+��b'����f�\q�yvG��%D�̬���J��*��]fF?�qIZt��J#�8w��GHe�:A"D&:��_+$)�����
7��O�{+�����QS�(��w�2uF��dԦ��;�����M�O�`����V�M�s�ܞK����9�̥��qތ���k0��3�c�� ��ߔ��P�A�v�q8z��O0 .ԏWg�Ce�w½�v)r���!�И����dR������sM��ۦ-/uxt���
�̮g�r��4� ��	��JEҧ��O]CJ<�Նg>r��M�&QUи�B�-7G��@�e� �����ʔ\�/eI@j�S��3�Y���ZC�����z&����X�Q�ʀ��HӦ�b����6�G��Bj��z��L������vߜ�*'�z5Ҕ~�ދ�Ĵh��_)i�.� m��D�R��d����0O-�(���ځB�����/|]�5��~�T����K�u��s��ް#�]gp�8�κ�4�jll藗��&؉5��e�Ex���p�U��@����#�F���08��x����H�r0Z��j5�lOC&���Q{�ÿg��{�Wޝ����ˤC���R��N�T��MF�D#���3!$�)a��$�ŀ,ut޺���lJ��Ѽ�x�&��|L%CIͬR�&��lU��֜��p�3e��Ӕ���t�!����6��f!hq���1	p�/��ڏl �o���<i�@b���hw��G�4�?z΀��ʛ�d����r��5���	Mt_2Q]Ӏ�q� p��ae�Eߕ<b��F(&����_";Ў�N+�<����F/�[{�l��Dʶ �O��$I�j�x03�!�v�����BXk1 )�]������w�ᗒ�xb�ol�6�_n,Ӆ*��lҦ�����-�~!&���nCDP��W-
��xH?�q�u�Ec����.�g�:Xa5�;���F=?eX�ڭ�!�{L]���F���O�+^qūd�t������jV��$�㦲c[���\�������p�~r�(�y��mG�Q�
^fcp�'|��ڔ	�c�5��/�)��&G���Q�����s�H���&j�����a�>��h��_[��D�D6�:p=C�]����|��p@��$����]�G��\�K )�}B�oGTw{w�4�o�v�"���p�����ɭ����'M�)��M�7�l�����2�Ul�6��u��eS�-�$(�����&�f��X�t�q/s8ͩ!A3|��.�NZ�i����>�������c�]�`�*F�)q�?6���ڳ����&x��o�O�]~N:���e�䒥�_a�ѵ&x1m>U,�;��u!{��1�.Lz�о��23����z���e�N�4���o>9%T4�̋�c��5�MJ��!�߹�����$4�g�z��/S��/���J S��L�{��M~��3��R���i{>��	�`�$�H3���|D��2#��uC�T)�o�-|: �I�'��8]��!뽎t��Ѡd̎[�?�^v�����ށ]��ű~�k�k�+xH�8C�������h��}L�zx��z.�J!�P�*��그;��L������!m��zf�X;�e��U�B�ECR� 5����x��-l2 ���u(Ŏ,p���?����,�ũ�cA��K��Hԃ|et#ڨ��Y;��D��"㒨-�>����e8�}C���.t" �w���?���Vgc�{q�㣃(�2��/g��N�s�(���=���5.A"S�(�J�a�MJ�=NQak� �r��=7��Q+L�X�%E��޹��Y�F��>��󟗖��US�����y��Z�Kx����Q�y��h�u�L���7�~���r �N�﮺eт8�v��<=W��ѴGE%��1�]��^�0���eeo So^��t,t�Mdl٥�����d�%WG��vXi_��n��;�V�r��`~
c�n�_W��:!r�S��_��t��{���4��rj4�?"X�S�;o@PE<=�5w;"�GR���F���K(yV��;��F,2���.&�����B��-'~�x�J'��TsHt�'�V0�P�hX�r��9G�[�����P'�2
��d���Le��BmҰ��٣��� �*q _v6�q���I4�KSԑם=�`��g��(�<�Z�)<�3K�ܳ9��I�]`�f�pɝ��o���j.wɡ�CN~4,���WkW�[#�6� #�9��Z������x{��D��	����UH{3;��z�0&�p�ǉ�u�+���a�	w*�o�K�5�%g{AEA����ָ���LX�����X5�Zm�����0�(z*�N�)��bqԵN1��8�-�P���H��v�M׬[}�gaqZ^J�w�T�����_Vg3&�	�f�� Wx[G���M��F��X/*��nuȋ�|��M�OZR���{
54;�u����8vh
r�\[��0J��?}���]���ܼ�jY�ZR��\^&3?M�Ĭ�v-�ۂGv��֋"$�]���j��̀<;�	i?E��kv-��n	C}Y�M�;�Ue�˩��?�Q+�Xt����p��L��Ҏ6q���"&l�V�z@� ��Mr%2���*�b�ڲ	F�KI�\]�H�wg�1���V�O�)�[����v��1�����@�'Lv�g>N�Y��=���T'A�.@X�P:���G 5{����oej�`1��V_$-x6a!��9M@�y��#^-��ۿ��Ѓ���ʗ��3v��)sgnI߄��Ģ��~�Z��~�3�5R��h1��l��_�C���b�Y�B��*:���x��Q��Cs�P�;�> �5~�x�a�]���t�h��i�e(X���N�S
,^��jR3[_�ۮ��DT~`ޫq%ӯ�#��{9Ғ�������D� >@ �C�%�4X�=��}�لܯ�U&}�&�M��$
�ffcr +��q�9ǘ�]�H���(�	2�U?[�+�[��@5z��B���M{���� ܪ��pV&�-#��9*�>6�^/H`L���qVȿ	Ya i�Z�޹C�����No��n�):�����_U��&��1}H�/M�B����K�x��*�"�d�Mf��f����x�[�B���5���ı�Q]� ����aewc�0��bCnػ�;�/>&?Q��-���q
�q�^�e�Y,�JƩ�H(��7�DZqf wAߞ�l��~{�^���--/��1�1\u*�M��P�����
�ec��ĵ.$Z�`!�k�pә�x�1�tc��Gma:�+$b2���ƌ�|����0z)�\��Xsd�?�m�����=bR{���Gr���� ��j�D��|� �#�]вʇe�R4:��]��7���	�ql9��'�1����a+��A����o!�O{��=�-���gGM4J3�U�)C�㱿�wڝ')��
	-�d �He[3�'��{wE�*k�F��Z@9�I+Թ�k��rF��e9��C���ȭ�*F�m鞡����F���CM4>�S�t_��J��0�&��8�s �2���CF����t�]Dl��ɻ��8\����K�vK��e�U߷~�d�`�W�z�@����ef3Ra��|^f`I>{yޘR�==��&���[�M�Mj!5C3#M�=���8*�g�|�㠂<%��c>���t�4��K��hsh��������b�O��{��G���(����A����C/�^R$#CD���א����.~��²T)�N�h��ē\ђG����Ldtv����F�2���+6E��QCjje~I����OHdٌ���*e嶇�ҁ[͞j�Ԓ��TVcF���р�_�Q����{>4D��\���?OѬ��n|Sw�L҄o5��'_��_��f-e/���"s�d���/��ǽYb���#)�,՝f�Y���+7y �<{��-�O1h�)��H5����]= ��R��Y�'�p4�/	��0ER\���`��{?�V�C5:$��[�lgA��L-��,K����#k6&_�&��˃zI5��d��=�n��{M�|�7>9��b���G��9c�Fݓ/�ZP۫���t�� �\��}�;�M���}��������W^�ȬZF��[����b����q0��R��<�*�l��M�a�Dx�npU��~��� �NZ�N;U��v����b��ÒW�7�gEm����K��gÑ����0�/E��ӑ;C��s�M7D|��� (���K���N�FETC$P��,r���XMc�ՁH�ӋI=�B����-E���%�����\T���� ��8|6.��/ �}�z8ע)a��"�V�Ytu;@�J|db��d��vv�p�����0��:<ɾ��F��}��%�&�]�P���/�W9Uߵ���M�%��W�KqX�J�?�5*�"Ef�Jr�q����b��~[(�Wҩ"3��p��%h��c2�YL�#w?7D��rxʗ�Z�Tǚ>�6?��[O_f�+"��tdE�gT$u;����*�r	w�
:,��Z�ˑ3�����ѣ��ѝ�Q��!���|�d��3R��∖���6��lU4�+m���s��� �}��H%o��-F��I]ѓ���<+au��/f�S<�M���̶����r1>1p0�Fc�E�\BgG�3epR���T"x]����
�>�a]����aS=/�)��������'ȇBd����i_`:Ó�7#�o���6ا�0����y�B��6�����Vj�ém�6��:�ѳR~m�}�g>7��g*���f��%�-i�j:e]��j�,�or_�2�������\&2R{��<OVX��� ��滒�ǰP�<��ōk� rr?7v��.�K։�(.ƙ/{�D���UU�W{���}��F��ӊB��GH�����=����T*D6H�(���J���������ιޙ���\��i���`�����J�H����v�U�Or��������+_ۣ��eBY����!��e6�|�c��W3�}%<�T�P2ư��֥:4������6dl8;����F������Ts���4�93p�Qh��J@f+#�[z:�b@�s�Ͽ���B�jF�Yg#���3�s�E�x|�_	�4Ӧ'#�㄄�>�-2�����M
�9�\l�}����6B[�_�^�)��&��'�sT� �u��9$߲R��xne�)�:�T��$�,�x�8'�G��#8����������_)�L�m	���E<W�Gz��+�U�+�Vt��xd�W�7:(�j�YN���݄{�ƅ��B������g{�	���P���K5_ؼً��A������R3*>��"�}�o���Ȟ�ʘ	��@�Ⱥ�&��p�z�7a��˭����r���Q���Кwa[����9ZQ)��\"Ѷ�Y"��m����q+	%�����2�}�ѥ8xj�q�Ѝ�^׫tŹ�k
J|�1HzH8��BNq��x�)�IJW��1oQ�7z,:�ќ�E<��B��ܾ8C�0���.��k6�)�D~LJ{*���FH�[��8�Y�������� ��J3ю\A^,s��H �t)�j�X�ѷc�A3��^%oA�n�쾲 .՞�o��e}�̓����xNc�:��=�a��"E�j�t�� �g��Ở��W�^Ln�
�A�2M�~��n�7E(��]���TCml��b}S!0��+��Quv��̑� H���0�;b9�0��~��#RϬϬ�<�aXHA�6�v�k����̘)�|}����}4��_�c���X�s�5��bPѤ+&�֜ºι�ͅ�}G�W��v.-�R�:�u��ѿ��A*], Z�?7��{�����F��}ƖB���|�￁ʆx烼<�֡��(i)S�/?�ƤO��1���9Ş�lC��v�ȿ�l�Cf��ԇ��c�N��i	� r��7u^r�5���x�LM�nsP�`X��Ui��&��셚���$��j�K��ٖ��֔�7�=#:�cm�CP�$i��ǘ��sD�*[
IGrt�E� *w���N�.a����B����&�1��Uk�����+�v�_oY��Lq�4��B��,N!�/��Ig�Ϩ�)����&�}� alҷ$D--��HIYD���x��(<{C�Dy=��ͺ�Ǯ���	��ʣn�bq��9��F=!Z���/"Lz��C`�iRk���n�u,�UPCW����T����7�M�7)}l5�1�Y��;���uA�)���i�:$��Թ�k~>q�	�Q��-8�a��Y�9n�3�}�s�&!���O/ygL�$�D�����=j���?7 TW��D̨����x�
��{�c��lW�o#�.�DƲ�~]?R+�c��A�}�0�u�X��o�a%�?�w�Ʊ8U�`�'�n��/f�񞾂<�03S+�(#��ۀ�v���r�8�����	����GV�eh�߅S����9�J����V9ѮE��zW��GX⣆)8Yj2q,�(���0����Iw`%u`OyDX,L�6�e�b��20��$k���(��g�_}s�E�	�,
�9l��y)M�a8�ػ����,��q,6Pk�&i���BǺ&���pwU�ZZ�aoh���!�����J��:��&8��T�)\8�G�!C��'���u��LO6�s�`#��� �ʓ��n�[�;L�I��*6u���LШw���^��ɣɊz���v1��g0�̗�dq���J�_D&�Å�Yυ�v��T�yTٵL�H�J�I��v��}�Ԝ�ძ��K�tP^��gдoݗŪ����ȍ7���[�N��w��u3�� �ަ������cm��O�@����]y�1@#߃]�vdK��	2�d��H�ZٝdJ1��t�T4굙�{�xC��M}V��Ee����A��]"&����y$w�|�i��0���u��~g;�TO����6��+մ�S�k~ة?�����Ng:ւS�>�T�ϰ�'0f���ׅ�i���(��;1e]�0U0>n�K����N����'D�1'Ѫi��'��s����"��R �+��uXh�+��a����L�n�|�8��޼�_6e����!BF�]6�	z�{E�<����G�%}�52$�m>�����������+3��=��Xn�(zJd�l�q�����Z�z(HOʇϻZ*��Tˎۆ�x�o���8QPK,VV�b���P(d������V����}'�k��YO;E�΋$�[�H�ځߑ��M�1�Sh��󲠄m���ٍ�\�()��61����Ф���h.�g�:'��X5=�-'���� �Å@T�C��W� ��%,�9o�s��J<T��w(Z�Q��gHD��w"F<���J�Gk�51\ӝF���>�f��N���M��5�&���ڷͽ���m"��lDU.��k��d'h�6�'m%1A����ʼ�H��X��b�f�Ǿ�CP�n5o�x6��Y���h��2���؋j�,�7~�ג��ؙ��`�C��d�dl�K��S�0k\&3������i���8E
w�;`�A�HIv(���O��꼍vwU%3��6bd� P�Hn��w!�����8/�*����Od�{�>Y#X�2�Qb�`Z�T2����V�~o���m;���a�# 7t�+eqX\BX�d:��by<?O�n+����`��a4e��V�9a�s�o[�c )��3�,�6:)�^7k���λ2��D��w�z������>/4�n��.\c��d�aY��"W|㹜4ea��a_�s�c�$��c�wb��l��.���r�\�Y�L���?x�3&���Ն��<�-�#���S_����,RX�]�
ʪ�r�ݎ�Tdg�k��(��%�����p�ҁ��BH��_g�AT`�-¯W�;I�&�6������q�hQ5x1$�ot�}{�`�sR��#���F��2Cs@�fm ȫ��Pp��'�aDc�m4xl���/L5P
R���@71�YH���2�]��`�e�{�{_��|ɿhok(ko���>k�*$)��!�UH#<Ջ@��=j~Y�eޏ�x��?1J$A��U=U���j��*��q���d4�#!�(P|9��Ʃ_���
��X&[�R�[U�#�O h����Z�K�����!�e\[��Ĳ��+|���,�(8��9�5���`�HK	^jα	��B�H�5��a��+
�5K��fa ��x�5V ��Ϧ��s�ZAm�о����#m��n]�Q6�%|�Kv5P��Ozu���%$)�^��ܤ!á�U�)��u�W��	�E�������f]��pv#�T�I��( ��!�������W���Č���;HX�ʶ��U8��A����D4'��nÇQM���jpp�+hQ$&�ʋ������y"� 2yɁ{ ^�֦�m���7�9[�q6�N��%�;2X_�'��t�t0���5�c�*�S��z����7,Gqx��k/�	)�CD�g �A��d��%u��P�dN�2[���r��7'^�R�NQV���|3���P�
�k%�A,���y�}3�S���h������J�sڟ�g�y�a�!��C�6f�����,<�,��T��e	��hF����lS�=�����@�sR���)��0v�Ef�29�_]��|Ks��P��R�VV�!6���q!Ba1��.G�F�r�(�v}�$p��y�cهz�=R�����X��̕�`��F|H$�At�K�WPvI����16EV}I��$"�\�ß;45��1���E�^��lB�
��Q9����������-�Ɉ���S�Av�<�`ݞ2¹~�<�,�5��EGs�-T����> ��������!.��
߀��Ú��κ�xL�$�2،�7 ����]��S��G8��9t%��gh��I����0�$ �riG(��W.���	1NL����:�Y�SԉTe����5��*�If�i��P (�u��sQ�{��)��$F̼k��bz%�AW
�V ��;����<a]F�~�Cnr�xuR9��%�9��s�1�9�S��<Z� ��S65�@�6�h�=����W����y�~4�%���8}.o��Ad��
r�������<�ڏ�"�����K��\ȯ��ם^��+5_i�~�	Ȯeb㭽1��E��\�z��Qȇ�ÓB�ݚ�ʋ�&T�~�BH���_wI�8vAJ��՚k����۫!AC���RË����mK�;}v�Y�R��g����I7Ɛ��>���co��>����\�>K1I�k�����������T���\Zf=d��ʏ��+�H��SU��ᏝtX77]�z�����g�l�7g+xShk7�V�:��GDn��.�>��������ޑv]��X=UqZ<HeE@����1��F����ڥO�f����������g,C���$�XP��$�@��B���zP{dR�'}��q/�MD����MڅIn�:L���|*��}iP�Q��(�Q�i�������1�$�[^�4��^f��vQ7u�F�G�6�Q�lhDy�*䚯DpE�M��$X@��C�5F����Y��J�e�zD��j��f�^�B7#�JuvZ�OY8F���pB7�B/�s�R���m'Y����w yZhg%��GR��_q��U�����W?�\��Y��/����g��PuP��=��m�w͞Y������p�:)�)�j�d�<����'{�Ӂ��C)��[����A��>�{��p�-bMjbZ��^G��H�Ԅn=����X)������}x@��8ݖp���:��Үl�ZO_�hd�����l��5�`S����ey���dzpFKę��$,���zV�i~����'�2o҅�3���@��R$�@kH�vZpvJ��J��Eýb��5h����.nw0[��°St�.�#c��v�]H3��m����
��0F� �:l�e�A[��kl_w���>���lSy
���˹|G��m[�ndḜs��怍s��݈��j#�5C؛�rϾ�
Uf�I4Ik�VB�{�^�X 4��5�L�L�栅���2Ǽ� �hN�ܰ�.p�?��q{s�wh�ʀ����oǶ��I4��=� ��2���i/�To�������5���͘�>@F`Y���q�J#/G}6�)O��zR/��%X��Fh.�j��J׮d9ss-q�3j���m��N����n�н2�����}�YW�QfA��.\�
�8qbКx�x�Ce��PtK�w��0�.P��MO(�g��>-t�%���Yx~�~,�?��^�p����p��0�[+��k|_�\7��-���m	D���#0�����Z�s��Q)��L_��klH%r�1nDs��S� �Qr���!z;*:[+N&�$f�M��q`f��ڻgAѷ͎	_�~9x�,d���c�Y/5�Z�kX�����Gu�o��l�q�B������k��G�j/U����ؽ���
V:aEڂ�j���{F��MN_�K�� �T�3 ��!j׳����e�9��C@:,
x:�D�v�D`��e׷=�����U�-ߤ���tYͰ��b����x���o��=���% �*dq���:�ct@t��\z��jAw#���,1r������U⎷'��.�S>Kh[b�'c,j!n\�d��-6�!|���+��NNk,0��ZU܋&X�oĞ]X�J����	�5RZ@���q�y�����N^ha1��t-�_��	<� �v�ґF��:#��]T��f��J��9�*4�W�_�2S�ƫ���� O!��᭗�W�gc�;,�e1BC��`�6ˍ(*Sy־t�L�y�+�<ff��w��Vq�[<�H�?���|Zd��Dz8��h���y?��,���"y؛���-̝��0���	4a;6|��*P�׆�ov�vB;��O,J&KD���+�1�a�������l1���G+P�N!���Dt0k�G�I�k���!%�k*^p���������^�=�
��}굢����:K#�t�`y^��B�*�_\�������!�T!�3�!	��M�u��g��3w8�s�-u%�E%��}Rmss+6O��8��h?}�����p�{�Q��7�T�Cn�1��Ҿ���@B��Ɉ�_U�e�x��K,W��*	�L
��+�Q��ǂ�_ Yt�4m�9���:L�˦���=�I�)����$~�{�nI(}>1�&O��渢�&�od&+"� ]��~Zd"���?!�R�ADT
�e@BH��^�7a�fG���GP�u��&6��W߫m]�7�>v�@�rD�(/YO�ę~��P���K��+�I"��{�0T��7�~�Y��ڜ����a�Dҏs43&(t��!Y�W�=�t���Yz� sK!b!l��a��f"
�q�'��Lr*F����l��̏��֝^��`�Y��%S��F���*�x�s��'W��C($�%?��9��!~K�Ax0�U�����![��NJ��Āl`hôgX;�{�˾��d�Ǘ�;٧�����qU����_~�T��笂����OL��t:�>o��)~\� Zo�����A��6:0�y�ǰ�cwK�d���!���#"�'�|(͜^#��ʚ9;��Ч>y��X.��L$���b�PQ+f/}�_�xxF���Qcc���m̔�n߯�;�`�=�?��f��0�!X�.��q�b��K�����4�oA�q,�����·���z��������ز_\����[�>��u��ܙ�������P�dX��gGةK��퓜��"L��g4[��{G�vЋ8�O�^0�C�L�w~<�05�K�Fc�m���j�)��l��=f�Oh�w�����:�����N�g@om��*#��=r��`{,�#@���kDDQ���,�q��W�2���U�e��?��*t� goÖu�e(D�+��^��N:G�`]�M��y���\ �,�=ƳH��ߊ���a)���`��p��\?�X�cǇN"����+�����c�(��J�Z�~� �I����o��C�B����|�r~� ��#�``�����@�r�Ym\�a��Z���T ���m��{ڽ�w��gN�nT�:o���!gY)��gV�f�&�;sݚ�a<���jQ9V̘}g\��4�&�{��i'�ཎ�8���طJ�+���+� ��$|��<�S�Q�����!y�łc��b3�y�րܓ�	
JD��]�JL�d�/7����e�Y]�[��(�O�Ϗ"��ņ�η	�`'a��B����X�'^���e`ڢ(���vU+�Ww��݄zn���S��Č���i䨈]ehV/[sޮד�ѫAP�x���0��.����)�~�zl�w{2�15Y�5G0,��]�e��^E[���?�&D�B�:��*	�[�Ɉ��~|p�3h�{����3�1�k7�E�*_"�	��`<����N�\
J%�t��ח�A��uv��/����:�l�A0��!�.��c �τ�KCܯ�La�ߝY���q��{�ks�B-�[��\�J;��"�E+���F�>||K�g
�G�����uvД�.�����q�B������Le�3��2�fP��=��j4��l��bJ�pw7b�-Ψ�e7�����~���-l9�����4�����"ϭp������Xx�c1}�G),�V��/R��?��&և���Wz-=˕q�������~���q
�վVh	�R��0ps���<K�Wo�^�ψG^biu�6>�l>�zWY¬����~�]&�S�9��!�x�^^EM���Ca���;QvF�-��_Bm�8�ZI|��ܑ[V*�@��)�,%?��e�q��'W��tD�%́Q�jYHf�R>E�	L0��<����^�Ee�Q:��p5���瘊�!|ęe��+(��qD7�������f`otV#�P]�n�f���b-���i�A�[R`e��__=��E�A9�GT\<�m�&�+��ް��
^>=��Vx�}P��E�L˯�]���L��q�F�L��V���
�>�1@9��?��Q�+�{�+��r����pY'�G���߸��b:C�=#�H{`���gi-=���U��yU�ǆ�$�����M��j�G�R�Z�R�';�"�X��``W��"����-)�N�)���]��������8:�&ް}�>s����֣	EFt!2�(���*PZ����X�\�M�ͤe,��clͻ:l]�(���9s&H��ʋ7'8�����XEF#( 8��g�1n�/c�S���?x��©׳䄂
� 5^Cց~;?M̑�&q���Zg�=��|飩��#f���,w�"�f�x�
p���=�O��Q_%M��u�d��*Y�=Wۇ��?�DV�(M��ub��-�|��=8��p� �o�V ��*�N����x,�~��-0��7����D�~�r$o��K�AǓ��n/!@�49�[C?��� �Á/��@�c6u�O�s1ԛ�'���%~�l^/tX�^0e	���<��N��׽�M�A�v#p>%�F%ѥʓI��챤�]-$WV��̖J�>������m�'�������������������4B��!#+o�1�����U�ߔ�����<V�u��W��p���(��te��D��[Bm�%���(�{P���GM���Ax�T��a2�.�
�"Š�i��1mM�g��FuAQh�
ӦQ�����/��`ıq���B�d(,�E~,����e3O�-�
p-��խ��ܶ�lK|���gn%��8�̟Tck)_U�x<hB��dDH��ݏ�8�RN�b��s�B�Q�6��_�b���q�6��� ���#�5�؜tL%?%V�QT¨����||U�;����x�De���W߅;�vW���Á�
R~�J�3k�
K��>��+�Â�q>4r��z�AP��lm3�e<"+/���,����}'(xcٯSu��+WWx]B������ǂ�5N��*�d�k��V๬�;v.�K�k4o�I��7��0�!.���;d����x良���Ί�-	��h��?��ϩ����>Vu��𕰬莅�m
�y�	n,ֹ��'�%
9���U�%9hq)�kN�V�����E��`��E�R��AL0�#��MJx9
�j���G��D�x���>��E�����+t�a$�@���(<R�fU)�:eM��!S�#��$Qx0����0�=�,J�����&-�̱�N'f쥠d�2� �z,<��r�
�)2'��(\I�>f3Z7ˎ39R4�{N���i�����̞�=j�&�Vd_����g�7���u � �X��� YE"S3���)��w|3tΖ�\0��e�fg��9gȜ��Q3{�ǻ�Ƌ%��,��oVkeCM|�`�K�V8�%�cK��}v�X[?�m�oB�U�&��G��0��i���iV4�jf(���,u_4���\�;������������׍�;mמn��F/�|u��$�.�t�3N<��{��B�Y�	>l=��;~)����F��+;	���Y�u���������F�qk�*�p3H����n�>��v�=2��~K���#�$��Q����0$B:�T����/�T�XN�Y7�/�M�GsهR��Z�)�O��H�_l_��<\~��G��qq.�PȦ�29�e�5䔭}m �*�W��Y̹_b��� �j�3�\jA2;굑ؓ�Q��݈��TݙW�R�C�ҕ��녝MT�E�J�Y'����R�C9*Ij��Y�P97���l2�Ԫ	�j���|F�cf��N��^�,
�t�]��i1j�<b�k�6������>�#�1;�p>�&Ǚ]Ne�y��8�ʹ*��Z�#a���8lޠ/۷�@+1 ��W����}�8t���[��()RDv��k���hFؒ���?�t���Ji�fI\
T]7��^b������_?���غH��z��"�u�#�,�$�1��_�Olh�MЈB�5^τL�����Oi伆
�݃Mљ��Qbk��S��>>{���%ǂ/�3�=�\Y����d�z�
�r����W��<���2���	�9ًQw�A",e�f6`"2��w.��:|�i������l:.���ߧ�pb/!a���ՠ:c+���	���2�J���=��i/��i3�q& v��DH�d��}G1㓂9P��,�Z%T�z}3m�.����ɦUjcڌ02��*E�S�U;g���7NF��)h��o�m�w���`��S9���5�~�����Q��1t��֭ &��Oc)���������}�@��uvT��|�^v��\�JԸ�*�x>_�czO2c{��&���cg�&�_<�,o_�E���۔{��M�@џ��IxJ��A��"]�-�
�S��8Cz��x�5
N�֮&/%�;�u���OP8-�wi����0��N�-�J�ӂ.���uY\�+��1o�d���܍qAK��8D׻��-AT@�f"7��j���*6◒�V�:�3�a�#���w�ನ[�i>�c�BT�Q�6:���o��紬�^�,�S-a���N�5V5�昽VRn����H_%�w���Hڰ�e��dU����?w&l���R��|�w03���6�6.4�j ���,�R^g,�L�5�������	"�ƚ���0������l+Mb�bP0�XQ]-��P�gY׉���;���rvG5��'qbh���%*kT���\�@$�F͑��O�*^H�o���+��QFv},�k�.�����p��yB���SD��]w���b�F7$��l�V^#T�OA�x�W�U�z������ ^��ҩy�a�������\.���Q�5���2EP4g�n��b����))�a���L@yD�����
� :�|rK�}D��$ vDl�i�<���<ٓ%t#U�lu8�9�ϔ�l}��5�xt�(	����l2b� ��^��J%�rlD-u��%�P�}�Z��2�QL̆P���t�����T�t�A^���ǒV3���U���0�ϰޅy�cyph��͝�F�[aU�Ie���4�*�ϐ���Z���w�Z40Lj7ޗ�ؘԵ3Ch|��O�a��`���w�bٞ���1�5;�'�U��<���%f��^|U�����cY)4ȡq�ϔ�ANes�Bt������<^}@NA�E�H�ږ����W���J9��g�iY<�Im]4�*|:��j�d���gf�lb���u� {�5����&@r#���.7���0�h�劲��̬b�}(�!d�|Ř�=����$�2��~ ���=����?Ɠۅ+���7��Ě*!�c�/)��WXR%�K7l�z�(�1�MwS��MKrEg���/\Y����ձF}��6�=�q)�+��<?���TL<}�_2�im)�!E^M�Y�ۏE6"RK8�/Ƶ��G��ǬvjP�oH�.�a���*�'"��{0���fr�x�_,oy��-P�C�3k��Ή�|�-3x4� ��@_[��'^�����RS�9��"Tx���]�5� zN.I��f���B�&�xSZ���/i�[��F�Yy�G��B�u{)�<�F���s�
P��fr1rF]���x�A��)��T�f�?�5W�@ h��,C���m����ʅL�C4�����x)w���>*o�p+��p*�6>ryI�L�ߧ��8�ˎ9�]W�>�ƈ
�"���`�Xٌ���������;�z���]rg��"I�K>񖕈��!+ڛ�.��p��ɱU|9����!I�E[Q����l�{�d�)JQ����x��M>����[��֮z��0�2I%a^�� Ӭ�(0�r��V�Ӣ�9��k�8�d7*(-�Xjg��x��+��@1�<;Z�F�ជf�S7��|_%������D���[P\F�=��ݢ�Mp�[[��i6*��c��n�)!<����/�_��O�#���̊q+-%#^a���n4a��*������6���ə%PХ���"���T�'�>i;=���� ��*$b<^�8t@<�T�uX�'Z��s�[����5���]c��E9r~�W6V�⮾���#X�M������Yhc<�p��}ͤ
�S5�%3o�0@j&��$��MG�bXrE7<�N��~S�����;rsKhJ���Hr��%��Ů��^�NO�.��r�g8���B����T�d�RG��_�u0rϒ�R�R��"m��ݞ��!�t�:��1+F�۔^�m"LEHT�V�	��a�͞� x�D��p�f�o8#�