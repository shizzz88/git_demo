  --Example instantiation for system 'my_processor'
  my_processor_inst : my_processor
    port map(
      LCD_E_from_the_lcd_0 => LCD_E_from_the_lcd_0,
      LCD_RS_from_the_lcd_0 => LCD_RS_from_the_lcd_0,
      LCD_RW_from_the_lcd_0 => LCD_RW_from_the_lcd_0,
      LCD_data_to_and_from_the_lcd_0 => LCD_data_to_and_from_the_lcd_0,
      MOSI_from_the_spi_0 => MOSI_from_the_spi_0,
      SCLK_from_the_spi_0 => SCLK_from_the_spi_0,
      SS_n_from_the_spi_0 => SS_n_from_the_spi_0,
      bidir_port_to_and_from_the_porta => bidir_port_to_and_from_the_porta,
      MISO_to_the_spi_0 => MISO_to_the_spi_0,
      clk_0 => clk_0,
      in_port_to_the_button => in_port_to_the_button,
      reset_n => reset_n
    );


